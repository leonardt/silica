

module corebit_and (
  input in0,
  input in1,
  output out
);
  assign out = in0 & in1;

endmodule //corebit_and

module corebit_or (
  input in0,
  input in1,
  output out
);
  assign out = in0 | in1;

endmodule //corebit_or

module coreir_or #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 | in1;

endmodule //coreir_or

module coreir_and #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 & in1;

endmodule //coreir_and

module corebit_const #(parameter value=1) (
  output out
);
  assign out = value;

endmodule //corebit_const

module coreir_add #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 + in1;

endmodule //coreir_add

module coreir_eq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 == in1;

endmodule //coreir_eq

module corebit_mux (
  input in0,
  input in1,
  input sel,
  output out
);
  assign out = sel ? in1 : in0;

endmodule //corebit_mux

module coreir_reg #(parameter init=1, parameter width=1) (
  input clk,
  input [width-1:0] in,
  output [width-1:0] out
);
reg [width-1:0] outReg=init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;

endmodule //coreir_reg

module or_wrapped (
  input  I0,
  input  I1,
  output  O
);
  //Wire declarations for instance 'inst0' (Module corebit_or)
  wire  inst0_in0;
  wire  inst0_out;
  wire  inst0_in1;
  corebit_or inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0 = I0;
  assign inst0_in1 = I1;
  assign O = inst0_out;

endmodule //or_wrapped

module Add2 (
  input [1:0] I0,
  input [1:0] I1,
  output [1:0] O
);
  //Wire declarations for instance 'inst0' (Module coreir_add)
  wire [1:0] inst0_in0;
  wire [1:0] inst0_out;
  wire [1:0] inst0_in1;
  coreir_add #(.width(2)) inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0[1:0] = I0[1:0];
  assign inst0_in1[1:0] = I1[1:0];
  assign O[1:0] = inst0_out[1:0];

endmodule //Add2

module corebit_not (
  input in,
  output out
);
  assign out = ~in;

endmodule //corebit_not

module EQ2 (
  input [1:0] I0,
  input [1:0] I1,
  output  O
);
  //Wire declarations for instance 'inst0' (Module coreir_eq)
  wire [1:0] inst0_in0;
  wire  inst0_out;
  wire [1:0] inst0_in1;
  coreir_eq #(.width(2)) inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0[1:0] = I0[1:0];
  assign inst0_in1[1:0] = I1[1:0];
  assign O = inst0_out;

endmodule //EQ2

module Decode22 (
  input [1:0] I,
  output  O
);
  //Wire declarations for instance 'bit_const_GND' (Module corebit_const)
  wire  bit_const_GND_out;
  corebit_const #(.value(0)) bit_const_GND(
    .out(bit_const_GND_out)
  );

  //Wire declarations for instance 'bit_const_VCC' (Module corebit_const)
  wire  bit_const_VCC_out;
  corebit_const #(.value(1)) bit_const_VCC(
    .out(bit_const_VCC_out)
  );

  //Wire declarations for instance 'inst0' (Module EQ2)
  wire [1:0] inst0_I0;
  wire [1:0] inst0_I1;
  wire  inst0_O;
  EQ2 inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //All the connections
  assign inst0_I1[0] = bit_const_GND_out;
  assign inst0_I1[1] = bit_const_VCC_out;
  assign inst0_I0[1:0] = I[1:0];
  assign O = inst0_O;

endmodule //Decode22

module Decode32 (
  input [1:0] I,
  output  O
);
  //Wire declarations for instance 'bit_const_VCC' (Module corebit_const)
  wire  bit_const_VCC_out;
  corebit_const #(.value(1)) bit_const_VCC(
    .out(bit_const_VCC_out)
  );

  //Wire declarations for instance 'inst0' (Module EQ2)
  wire [1:0] inst0_I0;
  wire [1:0] inst0_I1;
  wire  inst0_O;
  EQ2 inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //All the connections
  assign inst0_I1[0] = bit_const_VCC_out;
  assign inst0_I1[1] = bit_const_VCC_out;
  assign inst0_I0[1:0] = I[1:0];
  assign O = inst0_O;

endmodule //Decode32

module Decode02 (
  input [1:0] I,
  output  O
);
  //Wire declarations for instance 'bit_const_GND' (Module corebit_const)
  wire  bit_const_GND_out;
  corebit_const #(.value(0)) bit_const_GND(
    .out(bit_const_GND_out)
  );

  //Wire declarations for instance 'inst0' (Module EQ2)
  wire [1:0] inst0_I0;
  wire [1:0] inst0_I1;
  wire  inst0_O;
  EQ2 inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //All the connections
  assign inst0_I1[0] = bit_const_GND_out;
  assign inst0_I1[1] = bit_const_GND_out;
  assign inst0_I0[1:0] = I[1:0];
  assign O = inst0_O;

endmodule //Decode02

module Decode12 (
  input [1:0] I,
  output  O
);
  //Wire declarations for instance 'bit_const_GND' (Module corebit_const)
  wire  bit_const_GND_out;
  corebit_const #(.value(0)) bit_const_GND(
    .out(bit_const_GND_out)
  );

  //Wire declarations for instance 'bit_const_VCC' (Module corebit_const)
  wire  bit_const_VCC_out;
  corebit_const #(.value(1)) bit_const_VCC(
    .out(bit_const_VCC_out)
  );

  //Wire declarations for instance 'inst0' (Module EQ2)
  wire [1:0] inst0_I0;
  wire [1:0] inst0_I1;
  wire  inst0_O;
  EQ2 inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //All the connections
  assign inst0_I1[1] = bit_const_GND_out;
  assign inst0_I1[0] = bit_const_VCC_out;
  assign inst0_I0[1:0] = I[1:0];
  assign O = inst0_O;

endmodule //Decode12

module Decoder2 (
  input [1:0] I,
  output [3:0] O
);
  //Wire declarations for instance 'inst0' (Module Decode02)
  wire [1:0] inst0_I;
  wire  inst0_O;
  Decode02 inst0(
    .I(inst0_I),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module Decode12)
  wire [1:0] inst1_I;
  wire  inst1_O;
  Decode12 inst1(
    .I(inst1_I),
    .O(inst1_O)
  );

  //Wire declarations for instance 'inst2' (Module Decode22)
  wire [1:0] inst2_I;
  wire  inst2_O;
  Decode22 inst2(
    .I(inst2_I),
    .O(inst2_O)
  );

  //Wire declarations for instance 'inst3' (Module Decode32)
  wire [1:0] inst3_I;
  wire  inst3_O;
  Decode32 inst3(
    .I(inst3_I),
    .O(inst3_O)
  );

  //All the connections
  assign inst0_I[1:0] = I[1:0];
  assign O[0] = inst0_O;
  assign inst1_I[1:0] = I[1:0];
  assign O[1] = inst1_O;
  assign inst2_I[1:0] = I[1:0];
  assign O[2] = inst2_O;
  assign inst3_I[1:0] = I[1:0];
  assign O[3] = inst3_O;

endmodule //Decoder2

module _Mux2 (
  input [1:0] I,
  output  O,
  input  S
);
  //Wire declarations for instance 'inst0' (Module corebit_mux)
  wire  inst0_in0;
  wire  inst0_out;
  wire  inst0_in1;
  wire  inst0_sel;
  corebit_mux inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out),
    .sel(inst0_sel)
  );

  //All the connections
  assign inst0_in0 = I[0];
  assign inst0_in1 = I[1];
  assign O = inst0_out;
  assign inst0_sel = S;

endmodule //_Mux2

module _Mux4 (
  input [3:0] I,
  output  O,
  input [1:0] S
);
  //Wire declarations for instance 'inst0' (Module _Mux2)
  wire [1:0] inst0_I;
  wire  inst0_S;
  wire  inst0_O;
  _Mux2 inst0(
    .I(inst0_I),
    .O(inst0_O),
    .S(inst0_S)
  );

  //Wire declarations for instance 'inst1' (Module _Mux2)
  wire [1:0] inst1_I;
  wire  inst1_S;
  wire  inst1_O;
  _Mux2 inst1(
    .I(inst1_I),
    .O(inst1_O),
    .S(inst1_S)
  );

  //Wire declarations for instance 'inst2' (Module _Mux2)
  wire [1:0] inst2_I;
  wire  inst2_S;
  wire  inst2_O;
  _Mux2 inst2(
    .I(inst2_I),
    .O(inst2_O),
    .S(inst2_S)
  );

  //All the connections
  assign inst2_I[0] = inst0_O;
  assign inst0_S = S[0];
  assign inst2_I[1] = inst1_O;
  assign inst1_S = S[0];
  assign O = inst2_O;
  assign inst2_S = S[1];
  assign inst0_I[0] = I[0];
  assign inst0_I[1] = I[1];
  assign inst1_I[0] = I[2];
  assign inst1_I[1] = I[3];

endmodule //_Mux4

module Mux2x4 (
  input [3:0] I0,
  input [3:0] I1,
  output [3:0] O,
  input  S
);
  //Wire declarations for instance 'inst0' (Module _Mux2)
  wire [1:0] inst0_I;
  wire  inst0_S;
  wire  inst0_O;
  _Mux2 inst0(
    .I(inst0_I),
    .O(inst0_O),
    .S(inst0_S)
  );

  //Wire declarations for instance 'inst1' (Module _Mux2)
  wire [1:0] inst1_I;
  wire  inst1_S;
  wire  inst1_O;
  _Mux2 inst1(
    .I(inst1_I),
    .O(inst1_O),
    .S(inst1_S)
  );

  //Wire declarations for instance 'inst2' (Module _Mux2)
  wire [1:0] inst2_I;
  wire  inst2_S;
  wire  inst2_O;
  _Mux2 inst2(
    .I(inst2_I),
    .O(inst2_O),
    .S(inst2_S)
  );

  //Wire declarations for instance 'inst3' (Module _Mux2)
  wire [1:0] inst3_I;
  wire  inst3_S;
  wire  inst3_O;
  _Mux2 inst3(
    .I(inst3_I),
    .O(inst3_O),
    .S(inst3_S)
  );

  //All the connections
  assign O[0] = inst0_O;
  assign inst0_S = S;
  assign O[1] = inst1_O;
  assign inst1_S = S;
  assign O[2] = inst2_O;
  assign inst2_S = S;
  assign O[3] = inst3_O;
  assign inst3_S = S;
  assign inst0_I[0] = I0[0];
  assign inst0_I[1] = I1[0];
  assign inst1_I[0] = I0[1];
  assign inst1_I[1] = I1[1];
  assign inst2_I[0] = I0[2];
  assign inst2_I[1] = I1[2];
  assign inst3_I[0] = I0[3];
  assign inst3_I[1] = I1[3];

endmodule //Mux2x4

module Mux4x4 (
  input [3:0] I0,
  input [3:0] I1,
  input [3:0] I2,
  input [3:0] I3,
  output [3:0] O,
  input [1:0] S
);
  //Wire declarations for instance 'inst0' (Module _Mux4)
  wire [3:0] inst0_I;
  wire [1:0] inst0_S;
  wire  inst0_O;
  _Mux4 inst0(
    .I(inst0_I),
    .O(inst0_O),
    .S(inst0_S)
  );

  //Wire declarations for instance 'inst1' (Module _Mux4)
  wire [3:0] inst1_I;
  wire [1:0] inst1_S;
  wire  inst1_O;
  _Mux4 inst1(
    .I(inst1_I),
    .O(inst1_O),
    .S(inst1_S)
  );

  //Wire declarations for instance 'inst2' (Module _Mux4)
  wire [3:0] inst2_I;
  wire [1:0] inst2_S;
  wire  inst2_O;
  _Mux4 inst2(
    .I(inst2_I),
    .O(inst2_O),
    .S(inst2_S)
  );

  //Wire declarations for instance 'inst3' (Module _Mux4)
  wire [3:0] inst3_I;
  wire [1:0] inst3_S;
  wire  inst3_O;
  _Mux4 inst3(
    .I(inst3_I),
    .O(inst3_O),
    .S(inst3_S)
  );

  //All the connections
  assign O[0] = inst0_O;
  assign inst0_S[1:0] = S[1:0];
  assign O[1] = inst1_O;
  assign inst1_S[1:0] = S[1:0];
  assign O[2] = inst2_O;
  assign inst2_S[1:0] = S[1:0];
  assign O[3] = inst3_O;
  assign inst3_S[1:0] = S[1:0];
  assign inst0_I[0] = I0[0];
  assign inst0_I[1] = I1[0];
  assign inst0_I[2] = I2[0];
  assign inst0_I[3] = I3[0];
  assign inst1_I[0] = I0[1];
  assign inst1_I[1] = I1[1];
  assign inst1_I[2] = I2[1];
  assign inst1_I[3] = I3[1];
  assign inst2_I[0] = I0[2];
  assign inst2_I[1] = I1[2];
  assign inst2_I[2] = I2[2];
  assign inst2_I[3] = I3[2];
  assign inst3_I[0] = I0[3];
  assign inst3_I[1] = I1[3];
  assign inst3_I[2] = I2[3];
  assign inst3_I[3] = I3[3];

endmodule //Mux4x4

module reg_U1 #(parameter init=1) (
  input  clk,
  input [0:0] in,
  output [0:0] out
);
  //Wire declarations for instance 'reg0' (Module coreir_reg)
  wire  reg0_clk;
  wire [0:0] reg0_in;
  wire [0:0] reg0_out;
  coreir_reg #(.init(init),.width(1)) reg0(
    .clk(reg0_clk),
    .in(reg0_in),
    .out(reg0_out)
  );

  //All the connections
  assign reg0_clk = clk;
  assign reg0_in[0:0] = in[0:0];
  assign out[0:0] = reg0_out[0:0];

endmodule //reg_U1

module DFF_init0_has_ceFalse_has_resetFalse (
  input  CLK,
  input  I,
  output  O
);
  //Wire declarations for instance 'inst0' (Module reg_U1)
  wire [0:0] inst0_in;
  wire  inst0_clk;
  wire [0:0] inst0_out;
  reg_U1 #(.init(1'd0)) inst0(
    .clk(inst0_clk),
    .in(inst0_in),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_clk = CLK;
  assign inst0_in[0] = I;
  assign O = inst0_out[0];

endmodule //DFF_init0_has_ceFalse_has_resetFalse

module Register2 (
  input  CLK,
  input [1:0] I,
  output [1:0] O
);
  //Wire declarations for instance 'inst0' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst0_CLK;
  wire  inst0_I;
  wire  inst0_O;
  DFF_init0_has_ceFalse_has_resetFalse inst0(
    .CLK(inst0_CLK),
    .I(inst0_I),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst1_CLK;
  wire  inst1_I;
  wire  inst1_O;
  DFF_init0_has_ceFalse_has_resetFalse inst1(
    .CLK(inst1_CLK),
    .I(inst1_I),
    .O(inst1_O)
  );

  //All the connections
  assign inst0_CLK = CLK;
  assign inst0_I = I[0];
  assign O[0] = inst0_O;
  assign inst1_CLK = CLK;
  assign inst1_I = I[1];
  assign O[1] = inst1_O;

endmodule //Register2

module DFF_init1_has_ceFalse_has_resetFalse (
  input  CLK,
  input  I,
  output  O
);
  //Wire declarations for instance 'inst0' (Module reg_U1)
  wire [0:0] inst0_in;
  wire  inst0_clk;
  wire [0:0] inst0_out;
  reg_U1 #(.init(1'd1)) inst0(
    .clk(inst0_clk),
    .in(inst0_in),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_clk = CLK;
  assign inst0_in[0] = I;
  assign O = inst0_out[0];

endmodule //DFF_init1_has_ceFalse_has_resetFalse

module Register2_0001 (
  input  CLK,
  input [1:0] I,
  output [1:0] O
);
  //Wire declarations for instance 'inst0' (Module DFF_init1_has_ceFalse_has_resetFalse)
  wire  inst0_CLK;
  wire  inst0_I;
  wire  inst0_O;
  DFF_init1_has_ceFalse_has_resetFalse inst0(
    .CLK(inst0_CLK),
    .I(inst0_I),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst1_CLK;
  wire  inst1_I;
  wire  inst1_O;
  DFF_init0_has_ceFalse_has_resetFalse inst1(
    .CLK(inst1_CLK),
    .I(inst1_I),
    .O(inst1_O)
  );

  //All the connections
  assign inst0_CLK = CLK;
  assign inst0_I = I[0];
  assign O[0] = inst0_O;
  assign inst1_CLK = CLK;
  assign inst1_I = I[1];
  assign O[1] = inst1_O;

endmodule //Register2_0001

module Register4 (
  input  CLK,
  input [3:0] I,
  output [3:0] O
);
  //Wire declarations for instance 'inst0' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst0_CLK;
  wire  inst0_I;
  wire  inst0_O;
  DFF_init0_has_ceFalse_has_resetFalse inst0(
    .CLK(inst0_CLK),
    .I(inst0_I),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst1_CLK;
  wire  inst1_I;
  wire  inst1_O;
  DFF_init0_has_ceFalse_has_resetFalse inst1(
    .CLK(inst1_CLK),
    .I(inst1_I),
    .O(inst1_O)
  );

  //Wire declarations for instance 'inst2' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst2_CLK;
  wire  inst2_I;
  wire  inst2_O;
  DFF_init0_has_ceFalse_has_resetFalse inst2(
    .CLK(inst2_CLK),
    .I(inst2_I),
    .O(inst2_O)
  );

  //Wire declarations for instance 'inst3' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  inst3_CLK;
  wire  inst3_I;
  wire  inst3_O;
  DFF_init0_has_ceFalse_has_resetFalse inst3(
    .CLK(inst3_CLK),
    .I(inst3_I),
    .O(inst3_O)
  );

  //All the connections
  assign inst0_CLK = CLK;
  assign inst0_I = I[0];
  assign O[0] = inst0_O;
  assign inst1_CLK = CLK;
  assign inst1_I = I[1];
  assign O[1] = inst1_O;
  assign inst2_CLK = CLK;
  assign inst2_I = I[2];
  assign O[2] = inst2_O;
  assign inst3_CLK = CLK;
  assign inst3_I = I[3];
  assign O[3] = inst3_O;

endmodule //Register4

module __silica_BufferFifo (
  input [7:0] I,
  output [7:0] O
);
  //All the connections
  assign O[7:0] = I[7:0];

endmodule //__silica_BufferFifo

module and2_wrapped (
  input [1:0] I0,
  input [1:0] I1,
  output [1:0] O
);
  //Wire declarations for instance 'inst0' (Module coreir_and)
  wire [1:0] inst0_in0;
  wire [1:0] inst0_out;
  wire [1:0] inst0_in1;
  coreir_and #(.width(2)) inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0[1:0] = I0[1:0];
  assign inst0_in1[1:0] = I1[1:0];
  assign O[1:0] = inst0_out[1:0];

endmodule //and2_wrapped

module and4_wrapped (
  input [3:0] I0,
  input [3:0] I1,
  output [3:0] O
);
  //Wire declarations for instance 'inst0' (Module coreir_and)
  wire [3:0] inst0_in0;
  wire [3:0] inst0_out;
  wire [3:0] inst0_in1;
  coreir_and #(.width(4)) inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0[3:0] = I0[3:0];
  assign inst0_in1[3:0] = I1[3:0];
  assign O[3:0] = inst0_out[3:0];

endmodule //and4_wrapped

module and_wrapped (
  input  I0,
  input  I1,
  output  O
);
  //Wire declarations for instance 'inst0' (Module corebit_and)
  wire  inst0_in0;
  wire  inst0_out;
  wire  inst0_in1;
  corebit_and inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0 = I0;
  assign inst0_in1 = I1;
  assign O = inst0_out;

endmodule //and_wrapped

module fold_and3None (
  input  I0,
  input  I1,
  input  I2,
  output  O
);
  //Wire declarations for instance 'inst0' (Module and_wrapped)
  wire  inst0_I0;
  wire  inst0_I1;
  wire  inst0_O;
  and_wrapped inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module and_wrapped)
  wire  inst1_I0;
  wire  inst1_I1;
  wire  inst1_O;
  and_wrapped inst1(
    .I0(inst1_I0),
    .I1(inst1_I1),
    .O(inst1_O)
  );

  //All the connections
  assign inst0_I0 = I0;
  assign inst0_I1 = I1;
  assign inst1_I0 = inst0_O;
  assign inst1_I1 = I2;
  assign O = inst1_O;

endmodule //fold_and3None

module fold_or8None (
  input  I0,
  input  I1,
  input  I2,
  input  I3,
  input  I4,
  input  I5,
  input  I6,
  input  I7,
  output  O
);
  //Wire declarations for instance 'inst0' (Module or_wrapped)
  wire  inst0_I0;
  wire  inst0_I1;
  wire  inst0_O;
  or_wrapped inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module or_wrapped)
  wire  inst1_I0;
  wire  inst1_I1;
  wire  inst1_O;
  or_wrapped inst1(
    .I0(inst1_I0),
    .I1(inst1_I1),
    .O(inst1_O)
  );

  //Wire declarations for instance 'inst2' (Module or_wrapped)
  wire  inst2_I0;
  wire  inst2_I1;
  wire  inst2_O;
  or_wrapped inst2(
    .I0(inst2_I0),
    .I1(inst2_I1),
    .O(inst2_O)
  );

  //Wire declarations for instance 'inst3' (Module or_wrapped)
  wire  inst3_I0;
  wire  inst3_I1;
  wire  inst3_O;
  or_wrapped inst3(
    .I0(inst3_I0),
    .I1(inst3_I1),
    .O(inst3_O)
  );

  //Wire declarations for instance 'inst4' (Module or_wrapped)
  wire  inst4_I0;
  wire  inst4_I1;
  wire  inst4_O;
  or_wrapped inst4(
    .I0(inst4_I0),
    .I1(inst4_I1),
    .O(inst4_O)
  );

  //Wire declarations for instance 'inst5' (Module or_wrapped)
  wire  inst5_I0;
  wire  inst5_I1;
  wire  inst5_O;
  or_wrapped inst5(
    .I0(inst5_I0),
    .I1(inst5_I1),
    .O(inst5_O)
  );

  //Wire declarations for instance 'inst6' (Module or_wrapped)
  wire  inst6_I0;
  wire  inst6_I1;
  wire  inst6_O;
  or_wrapped inst6(
    .I0(inst6_I0),
    .I1(inst6_I1),
    .O(inst6_O)
  );

  //All the connections
  assign inst0_I0 = I0;
  assign inst0_I1 = I1;
  assign inst1_I0 = inst0_O;
  assign inst1_I1 = I2;
  assign inst2_I0 = inst1_O;
  assign inst2_I1 = I3;
  assign inst3_I0 = inst2_O;
  assign inst3_I1 = I4;
  assign inst4_I0 = inst3_O;
  assign inst4_I1 = I5;
  assign inst5_I0 = inst4_O;
  assign inst5_I1 = I6;
  assign inst6_I0 = inst5_O;
  assign inst6_I1 = I7;
  assign O = inst6_O;

endmodule //fold_or8None

module or2_wrapped (
  input [1:0] I0,
  input [1:0] I1,
  output [1:0] O
);
  //Wire declarations for instance 'inst0' (Module coreir_or)
  wire [1:0] inst0_in0;
  wire [1:0] inst0_out;
  wire [1:0] inst0_in1;
  coreir_or #(.width(2)) inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0[1:0] = I0[1:0];
  assign inst0_in1[1:0] = I1[1:0];
  assign O[1:0] = inst0_out[1:0];

endmodule //or2_wrapped

module fold_or82 (
  input [1:0] I0,
  input [1:0] I1,
  input [1:0] I2,
  input [1:0] I3,
  input [1:0] I4,
  input [1:0] I5,
  input [1:0] I6,
  input [1:0] I7,
  output [1:0] O
);
  //Wire declarations for instance 'inst0' (Module or2_wrapped)
  wire [1:0] inst0_I0;
  wire [1:0] inst0_I1;
  wire [1:0] inst0_O;
  or2_wrapped inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module or2_wrapped)
  wire [1:0] inst1_I0;
  wire [1:0] inst1_I1;
  wire [1:0] inst1_O;
  or2_wrapped inst1(
    .I0(inst1_I0),
    .I1(inst1_I1),
    .O(inst1_O)
  );

  //Wire declarations for instance 'inst2' (Module or2_wrapped)
  wire [1:0] inst2_I0;
  wire [1:0] inst2_I1;
  wire [1:0] inst2_O;
  or2_wrapped inst2(
    .I0(inst2_I0),
    .I1(inst2_I1),
    .O(inst2_O)
  );

  //Wire declarations for instance 'inst3' (Module or2_wrapped)
  wire [1:0] inst3_I0;
  wire [1:0] inst3_I1;
  wire [1:0] inst3_O;
  or2_wrapped inst3(
    .I0(inst3_I0),
    .I1(inst3_I1),
    .O(inst3_O)
  );

  //Wire declarations for instance 'inst4' (Module or2_wrapped)
  wire [1:0] inst4_I0;
  wire [1:0] inst4_I1;
  wire [1:0] inst4_O;
  or2_wrapped inst4(
    .I0(inst4_I0),
    .I1(inst4_I1),
    .O(inst4_O)
  );

  //Wire declarations for instance 'inst5' (Module or2_wrapped)
  wire [1:0] inst5_I0;
  wire [1:0] inst5_I1;
  wire [1:0] inst5_O;
  or2_wrapped inst5(
    .I0(inst5_I0),
    .I1(inst5_I1),
    .O(inst5_O)
  );

  //Wire declarations for instance 'inst6' (Module or2_wrapped)
  wire [1:0] inst6_I0;
  wire [1:0] inst6_I1;
  wire [1:0] inst6_O;
  or2_wrapped inst6(
    .I0(inst6_I0),
    .I1(inst6_I1),
    .O(inst6_O)
  );

  //All the connections
  assign inst0_I0[1:0] = I0[1:0];
  assign inst0_I1[1:0] = I1[1:0];
  assign inst1_I0[1:0] = inst0_O[1:0];
  assign inst1_I1[1:0] = I2[1:0];
  assign inst2_I0[1:0] = inst1_O[1:0];
  assign inst2_I1[1:0] = I3[1:0];
  assign inst3_I0[1:0] = inst2_O[1:0];
  assign inst3_I1[1:0] = I4[1:0];
  assign inst4_I0[1:0] = inst3_O[1:0];
  assign inst4_I1[1:0] = I5[1:0];
  assign inst5_I0[1:0] = inst4_O[1:0];
  assign inst5_I1[1:0] = I6[1:0];
  assign inst6_I0[1:0] = inst5_O[1:0];
  assign inst6_I1[1:0] = I7[1:0];
  assign O[1:0] = inst6_O[1:0];

endmodule //fold_or82

module or4_wrapped (
  input [3:0] I0,
  input [3:0] I1,
  output [3:0] O
);
  //Wire declarations for instance 'inst0' (Module coreir_or)
  wire [3:0] inst0_in0;
  wire [3:0] inst0_out;
  wire [3:0] inst0_in1;
  coreir_or #(.width(4)) inst0(
    .in0(inst0_in0),
    .in1(inst0_in1),
    .out(inst0_out)
  );

  //All the connections
  assign inst0_in0[3:0] = I0[3:0];
  assign inst0_in1[3:0] = I1[3:0];
  assign O[3:0] = inst0_out[3:0];

endmodule //or4_wrapped

module fold_or84 (
  input [3:0] I0,
  input [3:0] I1,
  input [3:0] I2,
  input [3:0] I3,
  input [3:0] I4,
  input [3:0] I5,
  input [3:0] I6,
  input [3:0] I7,
  output [3:0] O
);
  //Wire declarations for instance 'inst0' (Module or4_wrapped)
  wire [3:0] inst0_I0;
  wire [3:0] inst0_I1;
  wire [3:0] inst0_O;
  or4_wrapped inst0(
    .I0(inst0_I0),
    .I1(inst0_I1),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module or4_wrapped)
  wire [3:0] inst1_I0;
  wire [3:0] inst1_I1;
  wire [3:0] inst1_O;
  or4_wrapped inst1(
    .I0(inst1_I0),
    .I1(inst1_I1),
    .O(inst1_O)
  );

  //Wire declarations for instance 'inst2' (Module or4_wrapped)
  wire [3:0] inst2_I0;
  wire [3:0] inst2_I1;
  wire [3:0] inst2_O;
  or4_wrapped inst2(
    .I0(inst2_I0),
    .I1(inst2_I1),
    .O(inst2_O)
  );

  //Wire declarations for instance 'inst3' (Module or4_wrapped)
  wire [3:0] inst3_I0;
  wire [3:0] inst3_I1;
  wire [3:0] inst3_O;
  or4_wrapped inst3(
    .I0(inst3_I0),
    .I1(inst3_I1),
    .O(inst3_O)
  );

  //Wire declarations for instance 'inst4' (Module or4_wrapped)
  wire [3:0] inst4_I0;
  wire [3:0] inst4_I1;
  wire [3:0] inst4_O;
  or4_wrapped inst4(
    .I0(inst4_I0),
    .I1(inst4_I1),
    .O(inst4_O)
  );

  //Wire declarations for instance 'inst5' (Module or4_wrapped)
  wire [3:0] inst5_I0;
  wire [3:0] inst5_I1;
  wire [3:0] inst5_O;
  or4_wrapped inst5(
    .I0(inst5_I0),
    .I1(inst5_I1),
    .O(inst5_O)
  );

  //Wire declarations for instance 'inst6' (Module or4_wrapped)
  wire [3:0] inst6_I0;
  wire [3:0] inst6_I1;
  wire [3:0] inst6_O;
  or4_wrapped inst6(
    .I0(inst6_I0),
    .I1(inst6_I1),
    .O(inst6_O)
  );

  //All the connections
  assign inst0_I0[3:0] = I0[3:0];
  assign inst0_I1[3:0] = I1[3:0];
  assign inst1_I0[3:0] = inst0_O[3:0];
  assign inst1_I1[3:0] = I2[3:0];
  assign inst2_I0[3:0] = inst1_O[3:0];
  assign inst2_I1[3:0] = I3[3:0];
  assign inst3_I0[3:0] = inst2_O[3:0];
  assign inst3_I1[3:0] = I4[3:0];
  assign inst4_I0[3:0] = inst3_O[3:0];
  assign inst4_I1[3:0] = I5[3:0];
  assign inst5_I0[3:0] = inst4_O[3:0];
  assign inst5_I1[3:0] = I6[3:0];
  assign inst6_I0[3:0] = inst5_O[3:0];
  assign inst6_I1[3:0] = I7[3:0];
  assign O[3:0] = inst6_O[3:0];

endmodule //fold_or84

module Fifo (
  input  CLK,
  output  empty,
  output  full,
  output [3:0] rdata,
  input  ren,
  input [3:0] wdata,
  input  wen
);
  //Wire declarations for instance 'bit_const_GND' (Module corebit_const)
  wire  bit_const_GND_out;
  corebit_const #(.value(0)) bit_const_GND(
    .out(bit_const_GND_out)
  );

  //Wire declarations for instance 'bit_const_VCC' (Module corebit_const)
  wire  bit_const_VCC_out;
  corebit_const #(.value(1)) bit_const_VCC(
    .out(bit_const_VCC_out)
  );

  //Wire declarations for instance 'inst0' (Module __silica_BufferFifo)
  wire [7:0] inst0_I;
  wire [7:0] inst0_O;
  __silica_BufferFifo inst0(
    .I(inst0_I),
    .O(inst0_O)
  );

  //Wire declarations for instance 'inst1' (Module Register2_0001)
  wire  inst1_CLK;
  wire [1:0] inst1_I;
  wire [1:0] inst1_O;
  Register2_0001 inst1(
    .CLK(inst1_CLK),
    .I(inst1_I),
    .O(inst1_O)
  );

  //Wire declarations for instance 'inst10' (Module and2_wrapped)
  wire [1:0] inst10_I0;
  wire [1:0] inst10_I1;
  wire [1:0] inst10_O;
  and2_wrapped inst10(
    .I0(inst10_I0),
    .I1(inst10_I1),
    .O(inst10_O)
  );

  //Wire declarations for instance 'inst100' (Module fold_or8None)
  wire  inst100_I0;
  wire  inst100_I3;
  wire  inst100_O;
  wire  inst100_I4;
  wire  inst100_I2;
  wire  inst100_I1;
  wire  inst100_I7;
  wire  inst100_I5;
  wire  inst100_I6;
  fold_or8None inst100(
    .I0(inst100_I0),
    .I1(inst100_I1),
    .I2(inst100_I2),
    .I3(inst100_I3),
    .I4(inst100_I4),
    .I5(inst100_I5),
    .I6(inst100_I6),
    .I7(inst100_I7),
    .O(inst100_O)
  );

  //Wire declarations for instance 'inst101' (Module and_wrapped)
  wire  inst101_I0;
  wire  inst101_I1;
  wire  inst101_O;
  and_wrapped inst101(
    .I0(inst101_I0),
    .I1(inst101_I1),
    .O(inst101_O)
  );

  //Wire declarations for instance 'inst102' (Module and_wrapped)
  wire  inst102_I0;
  wire  inst102_I1;
  wire  inst102_O;
  and_wrapped inst102(
    .I0(inst102_I0),
    .I1(inst102_I1),
    .O(inst102_O)
  );

  //Wire declarations for instance 'inst103' (Module and_wrapped)
  wire  inst103_I0;
  wire  inst103_I1;
  wire  inst103_O;
  and_wrapped inst103(
    .I0(inst103_I0),
    .I1(inst103_I1),
    .O(inst103_O)
  );

  //Wire declarations for instance 'inst104' (Module and_wrapped)
  wire  inst104_I0;
  wire  inst104_I1;
  wire  inst104_O;
  and_wrapped inst104(
    .I0(inst104_I0),
    .I1(inst104_I1),
    .O(inst104_O)
  );

  //Wire declarations for instance 'inst105' (Module and_wrapped)
  wire  inst105_I0;
  wire  inst105_I1;
  wire  inst105_O;
  and_wrapped inst105(
    .I0(inst105_I0),
    .I1(inst105_I1),
    .O(inst105_O)
  );

  //Wire declarations for instance 'inst106' (Module and_wrapped)
  wire  inst106_I0;
  wire  inst106_I1;
  wire  inst106_O;
  and_wrapped inst106(
    .I0(inst106_I0),
    .I1(inst106_I1),
    .O(inst106_O)
  );

  //Wire declarations for instance 'inst107' (Module and_wrapped)
  wire  inst107_I0;
  wire  inst107_I1;
  wire  inst107_O;
  and_wrapped inst107(
    .I0(inst107_I0),
    .I1(inst107_I1),
    .O(inst107_O)
  );

  //Wire declarations for instance 'inst108' (Module and_wrapped)
  wire  inst108_I0;
  wire  inst108_I1;
  wire  inst108_O;
  and_wrapped inst108(
    .I0(inst108_I0),
    .I1(inst108_I1),
    .O(inst108_O)
  );

  //Wire declarations for instance 'inst109' (Module fold_or84)
  wire [3:0] inst109_I0;
  wire [3:0] inst109_I3;
  wire [3:0] inst109_O;
  wire [3:0] inst109_I4;
  wire [3:0] inst109_I2;
  wire [3:0] inst109_I1;
  wire [3:0] inst109_I7;
  wire [3:0] inst109_I5;
  wire [3:0] inst109_I6;
  fold_or84 inst109(
    .I0(inst109_I0),
    .I1(inst109_I1),
    .I2(inst109_I2),
    .I3(inst109_I3),
    .I4(inst109_I4),
    .I5(inst109_I5),
    .I6(inst109_I6),
    .I7(inst109_I7),
    .O(inst109_O)
  );

  //Wire declarations for instance 'inst11' (Module Register4)
  wire  inst11_CLK;
  wire [3:0] inst11_I;
  wire [3:0] inst11_O;
  Register4 inst11(
    .CLK(inst11_CLK),
    .I(inst11_I),
    .O(inst11_O)
  );

  //Wire declarations for instance 'inst110' (Module and4_wrapped)
  wire [3:0] inst110_I0;
  wire [3:0] inst110_I1;
  wire [3:0] inst110_O;
  and4_wrapped inst110(
    .I0(inst110_I0),
    .I1(inst110_I1),
    .O(inst110_O)
  );

  //Wire declarations for instance 'inst111' (Module and4_wrapped)
  wire [3:0] inst111_I0;
  wire [3:0] inst111_I1;
  wire [3:0] inst111_O;
  and4_wrapped inst111(
    .I0(inst111_I0),
    .I1(inst111_I1),
    .O(inst111_O)
  );

  //Wire declarations for instance 'inst112' (Module and4_wrapped)
  wire [3:0] inst112_I0;
  wire [3:0] inst112_I1;
  wire [3:0] inst112_O;
  and4_wrapped inst112(
    .I0(inst112_I0),
    .I1(inst112_I1),
    .O(inst112_O)
  );

  //Wire declarations for instance 'inst113' (Module and4_wrapped)
  wire [3:0] inst113_I0;
  wire [3:0] inst113_I1;
  wire [3:0] inst113_O;
  and4_wrapped inst113(
    .I0(inst113_I0),
    .I1(inst113_I1),
    .O(inst113_O)
  );

  //Wire declarations for instance 'inst114' (Module and4_wrapped)
  wire [3:0] inst114_I0;
  wire [3:0] inst114_I1;
  wire [3:0] inst114_O;
  and4_wrapped inst114(
    .I0(inst114_I0),
    .I1(inst114_I1),
    .O(inst114_O)
  );

  //Wire declarations for instance 'inst115' (Module and4_wrapped)
  wire [3:0] inst115_I0;
  wire [3:0] inst115_I1;
  wire [3:0] inst115_O;
  and4_wrapped inst115(
    .I0(inst115_I0),
    .I1(inst115_I1),
    .O(inst115_O)
  );

  //Wire declarations for instance 'inst116' (Module and4_wrapped)
  wire [3:0] inst116_I0;
  wire [3:0] inst116_I1;
  wire [3:0] inst116_O;
  and4_wrapped inst116(
    .I0(inst116_I0),
    .I1(inst116_I1),
    .O(inst116_O)
  );

  //Wire declarations for instance 'inst117' (Module and4_wrapped)
  wire [3:0] inst117_I0;
  wire [3:0] inst117_I1;
  wire [3:0] inst117_O;
  and4_wrapped inst117(
    .I0(inst117_I0),
    .I1(inst117_I1),
    .O(inst117_O)
  );

  //Wire declarations for instance 'inst118' (Module corebit_not)
  wire  inst118_in;
  wire  inst118_out;
  corebit_not inst118(
    .in(inst118_in),
    .out(inst118_out)
  );

  //Wire declarations for instance 'inst119' (Module and_wrapped)
  wire  inst119_I0;
  wire  inst119_I1;
  wire  inst119_O;
  and_wrapped inst119(
    .I0(inst119_I0),
    .I1(inst119_I1),
    .O(inst119_O)
  );

  //Wire declarations for instance 'inst12' (Module Register4)
  wire  inst12_CLK;
  wire [3:0] inst12_I;
  wire [3:0] inst12_O;
  Register4 inst12(
    .CLK(inst12_CLK),
    .I(inst12_I),
    .O(inst12_O)
  );

  //Wire declarations for instance 'inst120' (Module Decoder2)
  wire [1:0] inst120_I;
  wire [3:0] inst120_O;
  Decoder2 inst120(
    .I(inst120_I),
    .O(inst120_O)
  );

  //Wire declarations for instance 'inst121' (Module Mux2x4)
  wire [3:0] inst121_I0;
  wire [3:0] inst121_I1;
  wire [3:0] inst121_O;
  wire  inst121_S;
  Mux2x4 inst121(
    .I0(inst121_I0),
    .I1(inst121_I1),
    .O(inst121_O),
    .S(inst121_S)
  );

  //Wire declarations for instance 'inst122' (Module Mux2x4)
  wire [3:0] inst122_I0;
  wire [3:0] inst122_I1;
  wire [3:0] inst122_O;
  wire  inst122_S;
  Mux2x4 inst122(
    .I0(inst122_I0),
    .I1(inst122_I1),
    .O(inst122_O),
    .S(inst122_S)
  );

  //Wire declarations for instance 'inst123' (Module Mux2x4)
  wire [3:0] inst123_I0;
  wire [3:0] inst123_I1;
  wire [3:0] inst123_O;
  wire  inst123_S;
  Mux2x4 inst123(
    .I0(inst123_I0),
    .I1(inst123_I1),
    .O(inst123_O),
    .S(inst123_S)
  );

  //Wire declarations for instance 'inst124' (Module Mux2x4)
  wire [3:0] inst124_I0;
  wire [3:0] inst124_I1;
  wire [3:0] inst124_O;
  wire  inst124_S;
  Mux2x4 inst124(
    .I0(inst124_I0),
    .I1(inst124_I1),
    .O(inst124_O),
    .S(inst124_S)
  );

  //Wire declarations for instance 'inst125' (Module Add2)
  wire [1:0] inst125_I0;
  wire [1:0] inst125_I1;
  wire [1:0] inst125_O;
  Add2 inst125(
    .I0(inst125_I0),
    .I1(inst125_I1),
    .O(inst125_O)
  );

  //Wire declarations for instance 'inst126' (Module EQ2)
  wire [1:0] inst126_I0;
  wire [1:0] inst126_I1;
  wire  inst126_O;
  EQ2 inst126(
    .I0(inst126_I0),
    .I1(inst126_I1),
    .O(inst126_O)
  );

  //Wire declarations for instance 'inst127' (Module Mux4x4)
  wire [3:0] inst127_I0;
  wire [3:0] inst127_I1;
  wire [3:0] inst127_I2;
  wire [3:0] inst127_I3;
  wire [3:0] inst127_O;
  wire [1:0] inst127_S;
  Mux4x4 inst127(
    .I0(inst127_I0),
    .I1(inst127_I1),
    .I2(inst127_I2),
    .I3(inst127_I3),
    .O(inst127_O),
    .S(inst127_S)
  );

  //Wire declarations for instance 'inst128' (Module corebit_not)
  wire  inst128_in;
  wire  inst128_out;
  corebit_not inst128(
    .in(inst128_in),
    .out(inst128_out)
  );

  //Wire declarations for instance 'inst129' (Module and_wrapped)
  wire  inst129_I0;
  wire  inst129_I1;
  wire  inst129_O;
  and_wrapped inst129(
    .I0(inst129_I0),
    .I1(inst129_I1),
    .O(inst129_O)
  );

  //Wire declarations for instance 'inst13' (Module Register4)
  wire  inst13_CLK;
  wire [3:0] inst13_I;
  wire [3:0] inst13_O;
  Register4 inst13(
    .CLK(inst13_CLK),
    .I(inst13_I),
    .O(inst13_O)
  );

  //Wire declarations for instance 'inst130' (Module Add2)
  wire [1:0] inst130_I0;
  wire [1:0] inst130_I1;
  wire [1:0] inst130_O;
  Add2 inst130(
    .I0(inst130_I0),
    .I1(inst130_I1),
    .O(inst130_O)
  );

  //Wire declarations for instance 'inst131' (Module EQ2)
  wire [1:0] inst131_I0;
  wire [1:0] inst131_I1;
  wire  inst131_O;
  EQ2 inst131(
    .I0(inst131_I0),
    .I1(inst131_I1),
    .O(inst131_O)
  );

  //Wire declarations for instance 'inst132' (Module fold_and3None)
  wire  inst132_I0;
  wire  inst132_I1;
  wire  inst132_I2;
  wire  inst132_O;
  fold_and3None inst132(
    .I0(inst132_I0),
    .I1(inst132_I1),
    .I2(inst132_I2),
    .O(inst132_O)
  );

  //Wire declarations for instance 'inst133' (Module corebit_not)
  wire  inst133_in;
  wire  inst133_out;
  corebit_not inst133(
    .in(inst133_in),
    .out(inst133_out)
  );

  //Wire declarations for instance 'inst134' (Module and_wrapped)
  wire  inst134_I0;
  wire  inst134_I1;
  wire  inst134_O;
  and_wrapped inst134(
    .I0(inst134_I0),
    .I1(inst134_I1),
    .O(inst134_O)
  );

  //Wire declarations for instance 'inst135' (Module Decoder2)
  wire [1:0] inst135_I;
  wire [3:0] inst135_O;
  Decoder2 inst135(
    .I(inst135_I),
    .O(inst135_O)
  );

  //Wire declarations for instance 'inst136' (Module Mux2x4)
  wire [3:0] inst136_I0;
  wire [3:0] inst136_I1;
  wire [3:0] inst136_O;
  wire  inst136_S;
  Mux2x4 inst136(
    .I0(inst136_I0),
    .I1(inst136_I1),
    .O(inst136_O),
    .S(inst136_S)
  );

  //Wire declarations for instance 'inst137' (Module Mux2x4)
  wire [3:0] inst137_I0;
  wire [3:0] inst137_I1;
  wire [3:0] inst137_O;
  wire  inst137_S;
  Mux2x4 inst137(
    .I0(inst137_I0),
    .I1(inst137_I1),
    .O(inst137_O),
    .S(inst137_S)
  );

  //Wire declarations for instance 'inst138' (Module Mux2x4)
  wire [3:0] inst138_I0;
  wire [3:0] inst138_I1;
  wire [3:0] inst138_O;
  wire  inst138_S;
  Mux2x4 inst138(
    .I0(inst138_I0),
    .I1(inst138_I1),
    .O(inst138_O),
    .S(inst138_S)
  );

  //Wire declarations for instance 'inst139' (Module Mux2x4)
  wire [3:0] inst139_I0;
  wire [3:0] inst139_I1;
  wire [3:0] inst139_O;
  wire  inst139_S;
  Mux2x4 inst139(
    .I0(inst139_I0),
    .I1(inst139_I1),
    .O(inst139_O),
    .S(inst139_S)
  );

  //Wire declarations for instance 'inst14' (Module Register4)
  wire  inst14_CLK;
  wire [3:0] inst14_I;
  wire [3:0] inst14_O;
  Register4 inst14(
    .CLK(inst14_CLK),
    .I(inst14_I),
    .O(inst14_O)
  );

  //Wire declarations for instance 'inst140' (Module Add2)
  wire [1:0] inst140_I0;
  wire [1:0] inst140_I1;
  wire [1:0] inst140_O;
  Add2 inst140(
    .I0(inst140_I0),
    .I1(inst140_I1),
    .O(inst140_O)
  );

  //Wire declarations for instance 'inst141' (Module EQ2)
  wire [1:0] inst141_I0;
  wire [1:0] inst141_I1;
  wire  inst141_O;
  EQ2 inst141(
    .I0(inst141_I0),
    .I1(inst141_I1),
    .O(inst141_O)
  );

  //Wire declarations for instance 'inst142' (Module Mux4x4)
  wire [3:0] inst142_I0;
  wire [3:0] inst142_I1;
  wire [3:0] inst142_I2;
  wire [3:0] inst142_I3;
  wire [3:0] inst142_O;
  wire [1:0] inst142_S;
  Mux4x4 inst142(
    .I0(inst142_I0),
    .I1(inst142_I1),
    .I2(inst142_I2),
    .I3(inst142_I3),
    .O(inst142_O),
    .S(inst142_S)
  );

  //Wire declarations for instance 'inst143' (Module corebit_not)
  wire  inst143_in;
  wire  inst143_out;
  corebit_not inst143(
    .in(inst143_in),
    .out(inst143_out)
  );

  //Wire declarations for instance 'inst144' (Module and_wrapped)
  wire  inst144_I0;
  wire  inst144_I1;
  wire  inst144_O;
  and_wrapped inst144(
    .I0(inst144_I0),
    .I1(inst144_I1),
    .O(inst144_O)
  );

  //Wire declarations for instance 'inst145' (Module corebit_not)
  wire  inst145_in;
  wire  inst145_out;
  corebit_not inst145(
    .in(inst145_in),
    .out(inst145_out)
  );

  //Wire declarations for instance 'inst146' (Module fold_and3None)
  wire  inst146_I0;
  wire  inst146_I1;
  wire  inst146_I2;
  wire  inst146_O;
  fold_and3None inst146(
    .I0(inst146_I0),
    .I1(inst146_I1),
    .I2(inst146_I2),
    .O(inst146_O)
  );

  //Wire declarations for instance 'inst147' (Module corebit_not)
  wire  inst147_in;
  wire  inst147_out;
  corebit_not inst147(
    .in(inst147_in),
    .out(inst147_out)
  );

  //Wire declarations for instance 'inst148' (Module and_wrapped)
  wire  inst148_I0;
  wire  inst148_I1;
  wire  inst148_O;
  and_wrapped inst148(
    .I0(inst148_I0),
    .I1(inst148_I1),
    .O(inst148_O)
  );

  //Wire declarations for instance 'inst149' (Module corebit_not)
  wire  inst149_in;
  wire  inst149_out;
  corebit_not inst149(
    .in(inst149_in),
    .out(inst149_out)
  );

  //Wire declarations for instance 'inst15' (Module fold_or84)
  wire [3:0] inst15_I0;
  wire [3:0] inst15_I3;
  wire [3:0] inst15_O;
  wire [3:0] inst15_I4;
  wire [3:0] inst15_I2;
  wire [3:0] inst15_I1;
  wire [3:0] inst15_I7;
  wire [3:0] inst15_I5;
  wire [3:0] inst15_I6;
  fold_or84 inst15(
    .I0(inst15_I0),
    .I1(inst15_I1),
    .I2(inst15_I2),
    .I3(inst15_I3),
    .I4(inst15_I4),
    .I5(inst15_I5),
    .I6(inst15_I6),
    .I7(inst15_I7),
    .O(inst15_O)
  );

  //Wire declarations for instance 'inst150' (Module Mux4x4)
  wire [3:0] inst150_I0;
  wire [3:0] inst150_I1;
  wire [3:0] inst150_I2;
  wire [3:0] inst150_I3;
  wire [3:0] inst150_O;
  wire [1:0] inst150_S;
  Mux4x4 inst150(
    .I0(inst150_I0),
    .I1(inst150_I1),
    .I2(inst150_I2),
    .I3(inst150_I3),
    .O(inst150_O),
    .S(inst150_S)
  );

  //Wire declarations for instance 'inst151' (Module corebit_not)
  wire  inst151_in;
  wire  inst151_out;
  corebit_not inst151(
    .in(inst151_in),
    .out(inst151_out)
  );

  //Wire declarations for instance 'inst152' (Module and_wrapped)
  wire  inst152_I0;
  wire  inst152_I1;
  wire  inst152_O;
  and_wrapped inst152(
    .I0(inst152_I0),
    .I1(inst152_I1),
    .O(inst152_O)
  );

  //Wire declarations for instance 'inst153' (Module Add2)
  wire [1:0] inst153_I0;
  wire [1:0] inst153_I1;
  wire [1:0] inst153_O;
  Add2 inst153(
    .I0(inst153_I0),
    .I1(inst153_I1),
    .O(inst153_O)
  );

  //Wire declarations for instance 'inst154' (Module EQ2)
  wire [1:0] inst154_I0;
  wire [1:0] inst154_I1;
  wire  inst154_O;
  EQ2 inst154(
    .I0(inst154_I0),
    .I1(inst154_I1),
    .O(inst154_O)
  );

  //Wire declarations for instance 'inst155' (Module fold_and3None)
  wire  inst155_I0;
  wire  inst155_I1;
  wire  inst155_I2;
  wire  inst155_O;
  fold_and3None inst155(
    .I0(inst155_I0),
    .I1(inst155_I1),
    .I2(inst155_I2),
    .O(inst155_O)
  );

  //Wire declarations for instance 'inst156' (Module corebit_not)
  wire  inst156_in;
  wire  inst156_out;
  corebit_not inst156(
    .in(inst156_in),
    .out(inst156_out)
  );

  //Wire declarations for instance 'inst157' (Module and_wrapped)
  wire  inst157_I0;
  wire  inst157_I1;
  wire  inst157_O;
  and_wrapped inst157(
    .I0(inst157_I0),
    .I1(inst157_I1),
    .O(inst157_O)
  );

  //Wire declarations for instance 'inst158' (Module corebit_not)
  wire  inst158_in;
  wire  inst158_out;
  corebit_not inst158(
    .in(inst158_in),
    .out(inst158_out)
  );

  //Wire declarations for instance 'inst159' (Module Mux4x4)
  wire [3:0] inst159_I0;
  wire [3:0] inst159_I1;
  wire [3:0] inst159_I2;
  wire [3:0] inst159_I3;
  wire [3:0] inst159_O;
  wire [1:0] inst159_S;
  Mux4x4 inst159(
    .I0(inst159_I0),
    .I1(inst159_I1),
    .I2(inst159_I2),
    .I3(inst159_I3),
    .O(inst159_O),
    .S(inst159_S)
  );

  //Wire declarations for instance 'inst16' (Module fold_or84)
  wire [3:0] inst16_I0;
  wire [3:0] inst16_I3;
  wire [3:0] inst16_O;
  wire [3:0] inst16_I4;
  wire [3:0] inst16_I2;
  wire [3:0] inst16_I1;
  wire [3:0] inst16_I7;
  wire [3:0] inst16_I5;
  wire [3:0] inst16_I6;
  fold_or84 inst16(
    .I0(inst16_I0),
    .I1(inst16_I1),
    .I2(inst16_I2),
    .I3(inst16_I3),
    .I4(inst16_I4),
    .I5(inst16_I5),
    .I6(inst16_I6),
    .I7(inst16_I7),
    .O(inst16_O)
  );

  //Wire declarations for instance 'inst160' (Module corebit_not)
  wire  inst160_in;
  wire  inst160_out;
  corebit_not inst160(
    .in(inst160_in),
    .out(inst160_out)
  );

  //Wire declarations for instance 'inst161' (Module and_wrapped)
  wire  inst161_I0;
  wire  inst161_I1;
  wire  inst161_O;
  and_wrapped inst161(
    .I0(inst161_I0),
    .I1(inst161_I1),
    .O(inst161_O)
  );

  //Wire declarations for instance 'inst162' (Module corebit_not)
  wire  inst162_in;
  wire  inst162_out;
  corebit_not inst162(
    .in(inst162_in),
    .out(inst162_out)
  );

  //Wire declarations for instance 'inst163' (Module fold_and3None)
  wire  inst163_I0;
  wire  inst163_I1;
  wire  inst163_I2;
  wire  inst163_O;
  fold_and3None inst163(
    .I0(inst163_I0),
    .I1(inst163_I1),
    .I2(inst163_I2),
    .O(inst163_O)
  );

  //Wire declarations for instance 'inst164' (Module corebit_not)
  wire  inst164_in;
  wire  inst164_out;
  corebit_not inst164(
    .in(inst164_in),
    .out(inst164_out)
  );

  //Wire declarations for instance 'inst165' (Module and_wrapped)
  wire  inst165_I0;
  wire  inst165_I1;
  wire  inst165_O;
  and_wrapped inst165(
    .I0(inst165_I0),
    .I1(inst165_I1),
    .O(inst165_O)
  );

  //Wire declarations for instance 'inst166' (Module Decoder2)
  wire [1:0] inst166_I;
  wire [3:0] inst166_O;
  Decoder2 inst166(
    .I(inst166_I),
    .O(inst166_O)
  );

  //Wire declarations for instance 'inst167' (Module Mux2x4)
  wire [3:0] inst167_I0;
  wire [3:0] inst167_I1;
  wire [3:0] inst167_O;
  wire  inst167_S;
  Mux2x4 inst167(
    .I0(inst167_I0),
    .I1(inst167_I1),
    .O(inst167_O),
    .S(inst167_S)
  );

  //Wire declarations for instance 'inst168' (Module Mux2x4)
  wire [3:0] inst168_I0;
  wire [3:0] inst168_I1;
  wire [3:0] inst168_O;
  wire  inst168_S;
  Mux2x4 inst168(
    .I0(inst168_I0),
    .I1(inst168_I1),
    .O(inst168_O),
    .S(inst168_S)
  );

  //Wire declarations for instance 'inst169' (Module Mux2x4)
  wire [3:0] inst169_I0;
  wire [3:0] inst169_I1;
  wire [3:0] inst169_O;
  wire  inst169_S;
  Mux2x4 inst169(
    .I0(inst169_I0),
    .I1(inst169_I1),
    .O(inst169_O),
    .S(inst169_S)
  );

  //Wire declarations for instance 'inst17' (Module fold_or84)
  wire [3:0] inst17_I0;
  wire [3:0] inst17_I3;
  wire [3:0] inst17_O;
  wire [3:0] inst17_I4;
  wire [3:0] inst17_I2;
  wire [3:0] inst17_I1;
  wire [3:0] inst17_I7;
  wire [3:0] inst17_I5;
  wire [3:0] inst17_I6;
  fold_or84 inst17(
    .I0(inst17_I0),
    .I1(inst17_I1),
    .I2(inst17_I2),
    .I3(inst17_I3),
    .I4(inst17_I4),
    .I5(inst17_I5),
    .I6(inst17_I6),
    .I7(inst17_I7),
    .O(inst17_O)
  );

  //Wire declarations for instance 'inst170' (Module Mux2x4)
  wire [3:0] inst170_I0;
  wire [3:0] inst170_I1;
  wire [3:0] inst170_O;
  wire  inst170_S;
  Mux2x4 inst170(
    .I0(inst170_I0),
    .I1(inst170_I1),
    .O(inst170_O),
    .S(inst170_S)
  );

  //Wire declarations for instance 'inst171' (Module Add2)
  wire [1:0] inst171_I0;
  wire [1:0] inst171_I1;
  wire [1:0] inst171_O;
  Add2 inst171(
    .I0(inst171_I0),
    .I1(inst171_I1),
    .O(inst171_O)
  );

  //Wire declarations for instance 'inst172' (Module EQ2)
  wire [1:0] inst172_I0;
  wire [1:0] inst172_I1;
  wire  inst172_O;
  EQ2 inst172(
    .I0(inst172_I0),
    .I1(inst172_I1),
    .O(inst172_O)
  );

  //Wire declarations for instance 'inst173' (Module Mux4x4)
  wire [3:0] inst173_I0;
  wire [3:0] inst173_I1;
  wire [3:0] inst173_I2;
  wire [3:0] inst173_I3;
  wire [3:0] inst173_O;
  wire [1:0] inst173_S;
  Mux4x4 inst173(
    .I0(inst173_I0),
    .I1(inst173_I1),
    .I2(inst173_I2),
    .I3(inst173_I3),
    .O(inst173_O),
    .S(inst173_S)
  );

  //Wire declarations for instance 'inst174' (Module corebit_not)
  wire  inst174_in;
  wire  inst174_out;
  corebit_not inst174(
    .in(inst174_in),
    .out(inst174_out)
  );

  //Wire declarations for instance 'inst175' (Module and_wrapped)
  wire  inst175_I0;
  wire  inst175_I1;
  wire  inst175_O;
  and_wrapped inst175(
    .I0(inst175_I0),
    .I1(inst175_I1),
    .O(inst175_O)
  );

  //Wire declarations for instance 'inst176' (Module Add2)
  wire [1:0] inst176_I0;
  wire [1:0] inst176_I1;
  wire [1:0] inst176_O;
  Add2 inst176(
    .I0(inst176_I0),
    .I1(inst176_I1),
    .O(inst176_O)
  );

  //Wire declarations for instance 'inst177' (Module EQ2)
  wire [1:0] inst177_I0;
  wire [1:0] inst177_I1;
  wire  inst177_O;
  EQ2 inst177(
    .I0(inst177_I0),
    .I1(inst177_I1),
    .O(inst177_O)
  );

  //Wire declarations for instance 'inst178' (Module fold_and3None)
  wire  inst178_I0;
  wire  inst178_I1;
  wire  inst178_I2;
  wire  inst178_O;
  fold_and3None inst178(
    .I0(inst178_I0),
    .I1(inst178_I1),
    .I2(inst178_I2),
    .O(inst178_O)
  );

  //Wire declarations for instance 'inst179' (Module corebit_not)
  wire  inst179_in;
  wire  inst179_out;
  corebit_not inst179(
    .in(inst179_in),
    .out(inst179_out)
  );

  //Wire declarations for instance 'inst18' (Module fold_or84)
  wire [3:0] inst18_I0;
  wire [3:0] inst18_I3;
  wire [3:0] inst18_O;
  wire [3:0] inst18_I4;
  wire [3:0] inst18_I2;
  wire [3:0] inst18_I1;
  wire [3:0] inst18_I7;
  wire [3:0] inst18_I5;
  wire [3:0] inst18_I6;
  fold_or84 inst18(
    .I0(inst18_I0),
    .I1(inst18_I1),
    .I2(inst18_I2),
    .I3(inst18_I3),
    .I4(inst18_I4),
    .I5(inst18_I5),
    .I6(inst18_I6),
    .I7(inst18_I7),
    .O(inst18_O)
  );

  //Wire declarations for instance 'inst180' (Module and_wrapped)
  wire  inst180_I0;
  wire  inst180_I1;
  wire  inst180_O;
  and_wrapped inst180(
    .I0(inst180_I0),
    .I1(inst180_I1),
    .O(inst180_O)
  );

  //Wire declarations for instance 'inst181' (Module Decoder2)
  wire [1:0] inst181_I;
  wire [3:0] inst181_O;
  Decoder2 inst181(
    .I(inst181_I),
    .O(inst181_O)
  );

  //Wire declarations for instance 'inst182' (Module Mux2x4)
  wire [3:0] inst182_I0;
  wire [3:0] inst182_I1;
  wire [3:0] inst182_O;
  wire  inst182_S;
  Mux2x4 inst182(
    .I0(inst182_I0),
    .I1(inst182_I1),
    .O(inst182_O),
    .S(inst182_S)
  );

  //Wire declarations for instance 'inst183' (Module Mux2x4)
  wire [3:0] inst183_I0;
  wire [3:0] inst183_I1;
  wire [3:0] inst183_O;
  wire  inst183_S;
  Mux2x4 inst183(
    .I0(inst183_I0),
    .I1(inst183_I1),
    .O(inst183_O),
    .S(inst183_S)
  );

  //Wire declarations for instance 'inst184' (Module Mux2x4)
  wire [3:0] inst184_I0;
  wire [3:0] inst184_I1;
  wire [3:0] inst184_O;
  wire  inst184_S;
  Mux2x4 inst184(
    .I0(inst184_I0),
    .I1(inst184_I1),
    .O(inst184_O),
    .S(inst184_S)
  );

  //Wire declarations for instance 'inst185' (Module Mux2x4)
  wire [3:0] inst185_I0;
  wire [3:0] inst185_I1;
  wire [3:0] inst185_O;
  wire  inst185_S;
  Mux2x4 inst185(
    .I0(inst185_I0),
    .I1(inst185_I1),
    .O(inst185_O),
    .S(inst185_S)
  );

  //Wire declarations for instance 'inst186' (Module Add2)
  wire [1:0] inst186_I0;
  wire [1:0] inst186_I1;
  wire [1:0] inst186_O;
  Add2 inst186(
    .I0(inst186_I0),
    .I1(inst186_I1),
    .O(inst186_O)
  );

  //Wire declarations for instance 'inst187' (Module EQ2)
  wire [1:0] inst187_I0;
  wire [1:0] inst187_I1;
  wire  inst187_O;
  EQ2 inst187(
    .I0(inst187_I0),
    .I1(inst187_I1),
    .O(inst187_O)
  );

  //Wire declarations for instance 'inst188' (Module Mux4x4)
  wire [3:0] inst188_I0;
  wire [3:0] inst188_I1;
  wire [3:0] inst188_I2;
  wire [3:0] inst188_I3;
  wire [3:0] inst188_O;
  wire [1:0] inst188_S;
  Mux4x4 inst188(
    .I0(inst188_I0),
    .I1(inst188_I1),
    .I2(inst188_I2),
    .I3(inst188_I3),
    .O(inst188_O),
    .S(inst188_S)
  );

  //Wire declarations for instance 'inst189' (Module corebit_not)
  wire  inst189_in;
  wire  inst189_out;
  corebit_not inst189(
    .in(inst189_in),
    .out(inst189_out)
  );

  //Wire declarations for instance 'inst19' (Module and4_wrapped)
  wire [3:0] inst19_I0;
  wire [3:0] inst19_I1;
  wire [3:0] inst19_O;
  and4_wrapped inst19(
    .I0(inst19_I0),
    .I1(inst19_I1),
    .O(inst19_O)
  );

  //Wire declarations for instance 'inst190' (Module and_wrapped)
  wire  inst190_I0;
  wire  inst190_I1;
  wire  inst190_O;
  and_wrapped inst190(
    .I0(inst190_I0),
    .I1(inst190_I1),
    .O(inst190_O)
  );

  //Wire declarations for instance 'inst191' (Module corebit_not)
  wire  inst191_in;
  wire  inst191_out;
  corebit_not inst191(
    .in(inst191_in),
    .out(inst191_out)
  );

  //Wire declarations for instance 'inst192' (Module fold_and3None)
  wire  inst192_I0;
  wire  inst192_I1;
  wire  inst192_I2;
  wire  inst192_O;
  fold_and3None inst192(
    .I0(inst192_I0),
    .I1(inst192_I1),
    .I2(inst192_I2),
    .O(inst192_O)
  );

  //Wire declarations for instance 'inst193' (Module corebit_not)
  wire  inst193_in;
  wire  inst193_out;
  corebit_not inst193(
    .in(inst193_in),
    .out(inst193_out)
  );

  //Wire declarations for instance 'inst194' (Module and_wrapped)
  wire  inst194_I0;
  wire  inst194_I1;
  wire  inst194_O;
  and_wrapped inst194(
    .I0(inst194_I0),
    .I1(inst194_I1),
    .O(inst194_O)
  );

  //Wire declarations for instance 'inst195' (Module corebit_not)
  wire  inst195_in;
  wire  inst195_out;
  corebit_not inst195(
    .in(inst195_in),
    .out(inst195_out)
  );

  //Wire declarations for instance 'inst196' (Module Mux4x4)
  wire [3:0] inst196_I0;
  wire [3:0] inst196_I1;
  wire [3:0] inst196_I2;
  wire [3:0] inst196_I3;
  wire [3:0] inst196_O;
  wire [1:0] inst196_S;
  Mux4x4 inst196(
    .I0(inst196_I0),
    .I1(inst196_I1),
    .I2(inst196_I2),
    .I3(inst196_I3),
    .O(inst196_O),
    .S(inst196_S)
  );

  //Wire declarations for instance 'inst197' (Module corebit_not)
  wire  inst197_in;
  wire  inst197_out;
  corebit_not inst197(
    .in(inst197_in),
    .out(inst197_out)
  );

  //Wire declarations for instance 'inst198' (Module and_wrapped)
  wire  inst198_I0;
  wire  inst198_I1;
  wire  inst198_O;
  and_wrapped inst198(
    .I0(inst198_I0),
    .I1(inst198_I1),
    .O(inst198_O)
  );

  //Wire declarations for instance 'inst199' (Module Add2)
  wire [1:0] inst199_I0;
  wire [1:0] inst199_I1;
  wire [1:0] inst199_O;
  Add2 inst199(
    .I0(inst199_I0),
    .I1(inst199_I1),
    .O(inst199_O)
  );

  //Wire declarations for instance 'inst2' (Module fold_or82)
  wire [1:0] inst2_I0;
  wire [1:0] inst2_I3;
  wire [1:0] inst2_O;
  wire [1:0] inst2_I4;
  wire [1:0] inst2_I2;
  wire [1:0] inst2_I1;
  wire [1:0] inst2_I7;
  wire [1:0] inst2_I5;
  wire [1:0] inst2_I6;
  fold_or82 inst2(
    .I0(inst2_I0),
    .I1(inst2_I1),
    .I2(inst2_I2),
    .I3(inst2_I3),
    .I4(inst2_I4),
    .I5(inst2_I5),
    .I6(inst2_I6),
    .I7(inst2_I7),
    .O(inst2_O)
  );

  //Wire declarations for instance 'inst20' (Module and4_wrapped)
  wire [3:0] inst20_I0;
  wire [3:0] inst20_I1;
  wire [3:0] inst20_O;
  and4_wrapped inst20(
    .I0(inst20_I0),
    .I1(inst20_I1),
    .O(inst20_O)
  );

  //Wire declarations for instance 'inst200' (Module EQ2)
  wire [1:0] inst200_I0;
  wire [1:0] inst200_I1;
  wire  inst200_O;
  EQ2 inst200(
    .I0(inst200_I0),
    .I1(inst200_I1),
    .O(inst200_O)
  );

  //Wire declarations for instance 'inst201' (Module fold_and3None)
  wire  inst201_I0;
  wire  inst201_I1;
  wire  inst201_I2;
  wire  inst201_O;
  fold_and3None inst201(
    .I0(inst201_I0),
    .I1(inst201_I1),
    .I2(inst201_I2),
    .O(inst201_O)
  );

  //Wire declarations for instance 'inst202' (Module corebit_not)
  wire  inst202_in;
  wire  inst202_out;
  corebit_not inst202(
    .in(inst202_in),
    .out(inst202_out)
  );

  //Wire declarations for instance 'inst203' (Module and_wrapped)
  wire  inst203_I0;
  wire  inst203_I1;
  wire  inst203_O;
  and_wrapped inst203(
    .I0(inst203_I0),
    .I1(inst203_I1),
    .O(inst203_O)
  );

  //Wire declarations for instance 'inst204' (Module corebit_not)
  wire  inst204_in;
  wire  inst204_out;
  corebit_not inst204(
    .in(inst204_in),
    .out(inst204_out)
  );

  //Wire declarations for instance 'inst205' (Module Mux4x4)
  wire [3:0] inst205_I0;
  wire [3:0] inst205_I1;
  wire [3:0] inst205_I2;
  wire [3:0] inst205_I3;
  wire [3:0] inst205_O;
  wire [1:0] inst205_S;
  Mux4x4 inst205(
    .I0(inst205_I0),
    .I1(inst205_I1),
    .I2(inst205_I2),
    .I3(inst205_I3),
    .O(inst205_O),
    .S(inst205_S)
  );

  //Wire declarations for instance 'inst206' (Module corebit_not)
  wire  inst206_in;
  wire  inst206_out;
  corebit_not inst206(
    .in(inst206_in),
    .out(inst206_out)
  );

  //Wire declarations for instance 'inst207' (Module and_wrapped)
  wire  inst207_I0;
  wire  inst207_I1;
  wire  inst207_O;
  and_wrapped inst207(
    .I0(inst207_I0),
    .I1(inst207_I1),
    .O(inst207_O)
  );

  //Wire declarations for instance 'inst208' (Module corebit_not)
  wire  inst208_in;
  wire  inst208_out;
  corebit_not inst208(
    .in(inst208_in),
    .out(inst208_out)
  );

  //Wire declarations for instance 'inst209' (Module fold_and3None)
  wire  inst209_I0;
  wire  inst209_I1;
  wire  inst209_I2;
  wire  inst209_O;
  fold_and3None inst209(
    .I0(inst209_I0),
    .I1(inst209_I1),
    .I2(inst209_I2),
    .O(inst209_O)
  );

  //Wire declarations for instance 'inst21' (Module and4_wrapped)
  wire [3:0] inst21_I0;
  wire [3:0] inst21_I1;
  wire [3:0] inst21_O;
  and4_wrapped inst21(
    .I0(inst21_I0),
    .I1(inst21_I1),
    .O(inst21_O)
  );

  //Wire declarations for instance 'inst22' (Module and4_wrapped)
  wire [3:0] inst22_I0;
  wire [3:0] inst22_I1;
  wire [3:0] inst22_O;
  and4_wrapped inst22(
    .I0(inst22_I0),
    .I1(inst22_I1),
    .O(inst22_O)
  );

  //Wire declarations for instance 'inst23' (Module and4_wrapped)
  wire [3:0] inst23_I0;
  wire [3:0] inst23_I1;
  wire [3:0] inst23_O;
  and4_wrapped inst23(
    .I0(inst23_I0),
    .I1(inst23_I1),
    .O(inst23_O)
  );

  //Wire declarations for instance 'inst24' (Module and4_wrapped)
  wire [3:0] inst24_I0;
  wire [3:0] inst24_I1;
  wire [3:0] inst24_O;
  and4_wrapped inst24(
    .I0(inst24_I0),
    .I1(inst24_I1),
    .O(inst24_O)
  );

  //Wire declarations for instance 'inst25' (Module and4_wrapped)
  wire [3:0] inst25_I0;
  wire [3:0] inst25_I1;
  wire [3:0] inst25_O;
  and4_wrapped inst25(
    .I0(inst25_I0),
    .I1(inst25_I1),
    .O(inst25_O)
  );

  //Wire declarations for instance 'inst26' (Module and4_wrapped)
  wire [3:0] inst26_I0;
  wire [3:0] inst26_I1;
  wire [3:0] inst26_O;
  and4_wrapped inst26(
    .I0(inst26_I0),
    .I1(inst26_I1),
    .O(inst26_O)
  );

  //Wire declarations for instance 'inst27' (Module and4_wrapped)
  wire [3:0] inst27_I0;
  wire [3:0] inst27_I1;
  wire [3:0] inst27_O;
  and4_wrapped inst27(
    .I0(inst27_I0),
    .I1(inst27_I1),
    .O(inst27_O)
  );

  //Wire declarations for instance 'inst28' (Module and4_wrapped)
  wire [3:0] inst28_I0;
  wire [3:0] inst28_I1;
  wire [3:0] inst28_O;
  and4_wrapped inst28(
    .I0(inst28_I0),
    .I1(inst28_I1),
    .O(inst28_O)
  );

  //Wire declarations for instance 'inst29' (Module and4_wrapped)
  wire [3:0] inst29_I0;
  wire [3:0] inst29_I1;
  wire [3:0] inst29_O;
  and4_wrapped inst29(
    .I0(inst29_I0),
    .I1(inst29_I1),
    .O(inst29_O)
  );

  //Wire declarations for instance 'inst3' (Module and2_wrapped)
  wire [1:0] inst3_I0;
  wire [1:0] inst3_I1;
  wire [1:0] inst3_O;
  and2_wrapped inst3(
    .I0(inst3_I0),
    .I1(inst3_I1),
    .O(inst3_O)
  );

  //Wire declarations for instance 'inst30' (Module and4_wrapped)
  wire [3:0] inst30_I0;
  wire [3:0] inst30_I1;
  wire [3:0] inst30_O;
  and4_wrapped inst30(
    .I0(inst30_I0),
    .I1(inst30_I1),
    .O(inst30_O)
  );

  //Wire declarations for instance 'inst31' (Module and4_wrapped)
  wire [3:0] inst31_I0;
  wire [3:0] inst31_I1;
  wire [3:0] inst31_O;
  and4_wrapped inst31(
    .I0(inst31_I0),
    .I1(inst31_I1),
    .O(inst31_O)
  );

  //Wire declarations for instance 'inst32' (Module and4_wrapped)
  wire [3:0] inst32_I0;
  wire [3:0] inst32_I1;
  wire [3:0] inst32_O;
  and4_wrapped inst32(
    .I0(inst32_I0),
    .I1(inst32_I1),
    .O(inst32_O)
  );

  //Wire declarations for instance 'inst33' (Module and4_wrapped)
  wire [3:0] inst33_I0;
  wire [3:0] inst33_I1;
  wire [3:0] inst33_O;
  and4_wrapped inst33(
    .I0(inst33_I0),
    .I1(inst33_I1),
    .O(inst33_O)
  );

  //Wire declarations for instance 'inst34' (Module and4_wrapped)
  wire [3:0] inst34_I0;
  wire [3:0] inst34_I1;
  wire [3:0] inst34_O;
  and4_wrapped inst34(
    .I0(inst34_I0),
    .I1(inst34_I1),
    .O(inst34_O)
  );

  //Wire declarations for instance 'inst35' (Module and4_wrapped)
  wire [3:0] inst35_I0;
  wire [3:0] inst35_I1;
  wire [3:0] inst35_O;
  and4_wrapped inst35(
    .I0(inst35_I0),
    .I1(inst35_I1),
    .O(inst35_O)
  );

  //Wire declarations for instance 'inst36' (Module and4_wrapped)
  wire [3:0] inst36_I0;
  wire [3:0] inst36_I1;
  wire [3:0] inst36_O;
  and4_wrapped inst36(
    .I0(inst36_I0),
    .I1(inst36_I1),
    .O(inst36_O)
  );

  //Wire declarations for instance 'inst37' (Module and4_wrapped)
  wire [3:0] inst37_I0;
  wire [3:0] inst37_I1;
  wire [3:0] inst37_O;
  and4_wrapped inst37(
    .I0(inst37_I0),
    .I1(inst37_I1),
    .O(inst37_O)
  );

  //Wire declarations for instance 'inst38' (Module and4_wrapped)
  wire [3:0] inst38_I0;
  wire [3:0] inst38_I1;
  wire [3:0] inst38_O;
  and4_wrapped inst38(
    .I0(inst38_I0),
    .I1(inst38_I1),
    .O(inst38_O)
  );

  //Wire declarations for instance 'inst39' (Module and4_wrapped)
  wire [3:0] inst39_I0;
  wire [3:0] inst39_I1;
  wire [3:0] inst39_O;
  and4_wrapped inst39(
    .I0(inst39_I0),
    .I1(inst39_I1),
    .O(inst39_O)
  );

  //Wire declarations for instance 'inst4' (Module and2_wrapped)
  wire [1:0] inst4_I0;
  wire [1:0] inst4_I1;
  wire [1:0] inst4_O;
  and2_wrapped inst4(
    .I0(inst4_I0),
    .I1(inst4_I1),
    .O(inst4_O)
  );

  //Wire declarations for instance 'inst40' (Module and4_wrapped)
  wire [3:0] inst40_I0;
  wire [3:0] inst40_I1;
  wire [3:0] inst40_O;
  and4_wrapped inst40(
    .I0(inst40_I0),
    .I1(inst40_I1),
    .O(inst40_O)
  );

  //Wire declarations for instance 'inst41' (Module and4_wrapped)
  wire [3:0] inst41_I0;
  wire [3:0] inst41_I1;
  wire [3:0] inst41_O;
  and4_wrapped inst41(
    .I0(inst41_I0),
    .I1(inst41_I1),
    .O(inst41_O)
  );

  //Wire declarations for instance 'inst42' (Module and4_wrapped)
  wire [3:0] inst42_I0;
  wire [3:0] inst42_I1;
  wire [3:0] inst42_O;
  and4_wrapped inst42(
    .I0(inst42_I0),
    .I1(inst42_I1),
    .O(inst42_O)
  );

  //Wire declarations for instance 'inst43' (Module and4_wrapped)
  wire [3:0] inst43_I0;
  wire [3:0] inst43_I1;
  wire [3:0] inst43_O;
  and4_wrapped inst43(
    .I0(inst43_I0),
    .I1(inst43_I1),
    .O(inst43_O)
  );

  //Wire declarations for instance 'inst44' (Module and4_wrapped)
  wire [3:0] inst44_I0;
  wire [3:0] inst44_I1;
  wire [3:0] inst44_O;
  and4_wrapped inst44(
    .I0(inst44_I0),
    .I1(inst44_I1),
    .O(inst44_O)
  );

  //Wire declarations for instance 'inst45' (Module and4_wrapped)
  wire [3:0] inst45_I0;
  wire [3:0] inst45_I1;
  wire [3:0] inst45_O;
  and4_wrapped inst45(
    .I0(inst45_I0),
    .I1(inst45_I1),
    .O(inst45_O)
  );

  //Wire declarations for instance 'inst46' (Module and4_wrapped)
  wire [3:0] inst46_I0;
  wire [3:0] inst46_I1;
  wire [3:0] inst46_O;
  and4_wrapped inst46(
    .I0(inst46_I0),
    .I1(inst46_I1),
    .O(inst46_O)
  );

  //Wire declarations for instance 'inst47' (Module and4_wrapped)
  wire [3:0] inst47_I0;
  wire [3:0] inst47_I1;
  wire [3:0] inst47_O;
  and4_wrapped inst47(
    .I0(inst47_I0),
    .I1(inst47_I1),
    .O(inst47_O)
  );

  //Wire declarations for instance 'inst48' (Module and4_wrapped)
  wire [3:0] inst48_I0;
  wire [3:0] inst48_I1;
  wire [3:0] inst48_O;
  and4_wrapped inst48(
    .I0(inst48_I0),
    .I1(inst48_I1),
    .O(inst48_O)
  );

  //Wire declarations for instance 'inst49' (Module and4_wrapped)
  wire [3:0] inst49_I0;
  wire [3:0] inst49_I1;
  wire [3:0] inst49_O;
  and4_wrapped inst49(
    .I0(inst49_I0),
    .I1(inst49_I1),
    .O(inst49_O)
  );

  //Wire declarations for instance 'inst5' (Module and2_wrapped)
  wire [1:0] inst5_I0;
  wire [1:0] inst5_I1;
  wire [1:0] inst5_O;
  and2_wrapped inst5(
    .I0(inst5_I0),
    .I1(inst5_I1),
    .O(inst5_O)
  );

  //Wire declarations for instance 'inst50' (Module and4_wrapped)
  wire [3:0] inst50_I0;
  wire [3:0] inst50_I1;
  wire [3:0] inst50_O;
  and4_wrapped inst50(
    .I0(inst50_I0),
    .I1(inst50_I1),
    .O(inst50_O)
  );

  //Wire declarations for instance 'inst51' (Module Register2)
  wire  inst51_CLK;
  wire [1:0] inst51_I;
  wire [1:0] inst51_O;
  Register2 inst51(
    .CLK(inst51_CLK),
    .I(inst51_I),
    .O(inst51_O)
  );

  //Wire declarations for instance 'inst52' (Module fold_or82)
  wire [1:0] inst52_I0;
  wire [1:0] inst52_I3;
  wire [1:0] inst52_O;
  wire [1:0] inst52_I4;
  wire [1:0] inst52_I2;
  wire [1:0] inst52_I1;
  wire [1:0] inst52_I7;
  wire [1:0] inst52_I5;
  wire [1:0] inst52_I6;
  fold_or82 inst52(
    .I0(inst52_I0),
    .I1(inst52_I1),
    .I2(inst52_I2),
    .I3(inst52_I3),
    .I4(inst52_I4),
    .I5(inst52_I5),
    .I6(inst52_I6),
    .I7(inst52_I7),
    .O(inst52_O)
  );

  //Wire declarations for instance 'inst53' (Module and2_wrapped)
  wire [1:0] inst53_I0;
  wire [1:0] inst53_I1;
  wire [1:0] inst53_O;
  and2_wrapped inst53(
    .I0(inst53_I0),
    .I1(inst53_I1),
    .O(inst53_O)
  );

  //Wire declarations for instance 'inst54' (Module and2_wrapped)
  wire [1:0] inst54_I0;
  wire [1:0] inst54_I1;
  wire [1:0] inst54_O;
  and2_wrapped inst54(
    .I0(inst54_I0),
    .I1(inst54_I1),
    .O(inst54_O)
  );

  //Wire declarations for instance 'inst55' (Module and2_wrapped)
  wire [1:0] inst55_I0;
  wire [1:0] inst55_I1;
  wire [1:0] inst55_O;
  and2_wrapped inst55(
    .I0(inst55_I0),
    .I1(inst55_I1),
    .O(inst55_O)
  );

  //Wire declarations for instance 'inst56' (Module and2_wrapped)
  wire [1:0] inst56_I0;
  wire [1:0] inst56_I1;
  wire [1:0] inst56_O;
  and2_wrapped inst56(
    .I0(inst56_I0),
    .I1(inst56_I1),
    .O(inst56_O)
  );

  //Wire declarations for instance 'inst57' (Module and2_wrapped)
  wire [1:0] inst57_I0;
  wire [1:0] inst57_I1;
  wire [1:0] inst57_O;
  and2_wrapped inst57(
    .I0(inst57_I0),
    .I1(inst57_I1),
    .O(inst57_O)
  );

  //Wire declarations for instance 'inst58' (Module and2_wrapped)
  wire [1:0] inst58_I0;
  wire [1:0] inst58_I1;
  wire [1:0] inst58_O;
  and2_wrapped inst58(
    .I0(inst58_I0),
    .I1(inst58_I1),
    .O(inst58_O)
  );

  //Wire declarations for instance 'inst59' (Module and2_wrapped)
  wire [1:0] inst59_I0;
  wire [1:0] inst59_I1;
  wire [1:0] inst59_O;
  and2_wrapped inst59(
    .I0(inst59_I0),
    .I1(inst59_I1),
    .O(inst59_O)
  );

  //Wire declarations for instance 'inst6' (Module and2_wrapped)
  wire [1:0] inst6_I0;
  wire [1:0] inst6_I1;
  wire [1:0] inst6_O;
  and2_wrapped inst6(
    .I0(inst6_I0),
    .I1(inst6_I1),
    .O(inst6_O)
  );

  //Wire declarations for instance 'inst60' (Module and2_wrapped)
  wire [1:0] inst60_I0;
  wire [1:0] inst60_I1;
  wire [1:0] inst60_O;
  and2_wrapped inst60(
    .I0(inst60_I0),
    .I1(inst60_I1),
    .O(inst60_O)
  );

  //Wire declarations for instance 'inst61' (Module Register2)
  wire  inst61_CLK;
  wire [1:0] inst61_I;
  wire [1:0] inst61_O;
  Register2 inst61(
    .CLK(inst61_CLK),
    .I(inst61_I),
    .O(inst61_O)
  );

  //Wire declarations for instance 'inst62' (Module fold_or82)
  wire [1:0] inst62_I0;
  wire [1:0] inst62_I3;
  wire [1:0] inst62_O;
  wire [1:0] inst62_I4;
  wire [1:0] inst62_I2;
  wire [1:0] inst62_I1;
  wire [1:0] inst62_I7;
  wire [1:0] inst62_I5;
  wire [1:0] inst62_I6;
  fold_or82 inst62(
    .I0(inst62_I0),
    .I1(inst62_I1),
    .I2(inst62_I2),
    .I3(inst62_I3),
    .I4(inst62_I4),
    .I5(inst62_I5),
    .I6(inst62_I6),
    .I7(inst62_I7),
    .O(inst62_O)
  );

  //Wire declarations for instance 'inst63' (Module and2_wrapped)
  wire [1:0] inst63_I0;
  wire [1:0] inst63_I1;
  wire [1:0] inst63_O;
  and2_wrapped inst63(
    .I0(inst63_I0),
    .I1(inst63_I1),
    .O(inst63_O)
  );

  //Wire declarations for instance 'inst64' (Module and2_wrapped)
  wire [1:0] inst64_I0;
  wire [1:0] inst64_I1;
  wire [1:0] inst64_O;
  and2_wrapped inst64(
    .I0(inst64_I0),
    .I1(inst64_I1),
    .O(inst64_O)
  );

  //Wire declarations for instance 'inst65' (Module and2_wrapped)
  wire [1:0] inst65_I0;
  wire [1:0] inst65_I1;
  wire [1:0] inst65_O;
  and2_wrapped inst65(
    .I0(inst65_I0),
    .I1(inst65_I1),
    .O(inst65_O)
  );

  //Wire declarations for instance 'inst66' (Module and2_wrapped)
  wire [1:0] inst66_I0;
  wire [1:0] inst66_I1;
  wire [1:0] inst66_O;
  and2_wrapped inst66(
    .I0(inst66_I0),
    .I1(inst66_I1),
    .O(inst66_O)
  );

  //Wire declarations for instance 'inst67' (Module and2_wrapped)
  wire [1:0] inst67_I0;
  wire [1:0] inst67_I1;
  wire [1:0] inst67_O;
  and2_wrapped inst67(
    .I0(inst67_I0),
    .I1(inst67_I1),
    .O(inst67_O)
  );

  //Wire declarations for instance 'inst68' (Module and2_wrapped)
  wire [1:0] inst68_I0;
  wire [1:0] inst68_I1;
  wire [1:0] inst68_O;
  and2_wrapped inst68(
    .I0(inst68_I0),
    .I1(inst68_I1),
    .O(inst68_O)
  );

  //Wire declarations for instance 'inst69' (Module and2_wrapped)
  wire [1:0] inst69_I0;
  wire [1:0] inst69_I1;
  wire [1:0] inst69_O;
  and2_wrapped inst69(
    .I0(inst69_I0),
    .I1(inst69_I1),
    .O(inst69_O)
  );

  //Wire declarations for instance 'inst7' (Module and2_wrapped)
  wire [1:0] inst7_I0;
  wire [1:0] inst7_I1;
  wire [1:0] inst7_O;
  and2_wrapped inst7(
    .I0(inst7_I0),
    .I1(inst7_I1),
    .O(inst7_O)
  );

  //Wire declarations for instance 'inst70' (Module and2_wrapped)
  wire [1:0] inst70_I0;
  wire [1:0] inst70_I1;
  wire [1:0] inst70_O;
  and2_wrapped inst70(
    .I0(inst70_I0),
    .I1(inst70_I1),
    .O(inst70_O)
  );

  //Wire declarations for instance 'inst72' (Module fold_or8None)
  wire  inst72_I0;
  wire  inst72_I3;
  wire  inst72_O;
  wire  inst72_I4;
  wire  inst72_I2;
  wire  inst72_I1;
  wire  inst72_I7;
  wire  inst72_I5;
  wire  inst72_I6;
  fold_or8None inst72(
    .I0(inst72_I0),
    .I1(inst72_I1),
    .I2(inst72_I2),
    .I3(inst72_I3),
    .I4(inst72_I4),
    .I5(inst72_I5),
    .I6(inst72_I6),
    .I7(inst72_I7),
    .O(inst72_O)
  );

  //Wire declarations for instance 'inst73' (Module and_wrapped)
  wire  inst73_I0;
  wire  inst73_I1;
  wire  inst73_O;
  and_wrapped inst73(
    .I0(inst73_I0),
    .I1(inst73_I1),
    .O(inst73_O)
  );

  //Wire declarations for instance 'inst74' (Module and_wrapped)
  wire  inst74_I0;
  wire  inst74_I1;
  wire  inst74_O;
  and_wrapped inst74(
    .I0(inst74_I0),
    .I1(inst74_I1),
    .O(inst74_O)
  );

  //Wire declarations for instance 'inst75' (Module and_wrapped)
  wire  inst75_I0;
  wire  inst75_I1;
  wire  inst75_O;
  and_wrapped inst75(
    .I0(inst75_I0),
    .I1(inst75_I1),
    .O(inst75_O)
  );

  //Wire declarations for instance 'inst76' (Module and_wrapped)
  wire  inst76_I0;
  wire  inst76_I1;
  wire  inst76_O;
  and_wrapped inst76(
    .I0(inst76_I0),
    .I1(inst76_I1),
    .O(inst76_O)
  );

  //Wire declarations for instance 'inst77' (Module and_wrapped)
  wire  inst77_I0;
  wire  inst77_I1;
  wire  inst77_O;
  and_wrapped inst77(
    .I0(inst77_I0),
    .I1(inst77_I1),
    .O(inst77_O)
  );

  //Wire declarations for instance 'inst78' (Module and_wrapped)
  wire  inst78_I0;
  wire  inst78_I1;
  wire  inst78_O;
  and_wrapped inst78(
    .I0(inst78_I0),
    .I1(inst78_I1),
    .O(inst78_O)
  );

  //Wire declarations for instance 'inst79' (Module and_wrapped)
  wire  inst79_I0;
  wire  inst79_I1;
  wire  inst79_O;
  and_wrapped inst79(
    .I0(inst79_I0),
    .I1(inst79_I1),
    .O(inst79_O)
  );

  //Wire declarations for instance 'inst8' (Module and2_wrapped)
  wire [1:0] inst8_I0;
  wire [1:0] inst8_I1;
  wire [1:0] inst8_O;
  and2_wrapped inst8(
    .I0(inst8_I0),
    .I1(inst8_I1),
    .O(inst8_O)
  );

  //Wire declarations for instance 'inst80' (Module and_wrapped)
  wire  inst80_I0;
  wire  inst80_I1;
  wire  inst80_O;
  and_wrapped inst80(
    .I0(inst80_I0),
    .I1(inst80_I1),
    .O(inst80_O)
  );

  //Wire declarations for instance 'inst82' (Module fold_or8None)
  wire  inst82_I0;
  wire  inst82_I3;
  wire  inst82_O;
  wire  inst82_I4;
  wire  inst82_I2;
  wire  inst82_I1;
  wire  inst82_I7;
  wire  inst82_I5;
  wire  inst82_I6;
  fold_or8None inst82(
    .I0(inst82_I0),
    .I1(inst82_I1),
    .I2(inst82_I2),
    .I3(inst82_I3),
    .I4(inst82_I4),
    .I5(inst82_I5),
    .I6(inst82_I6),
    .I7(inst82_I7),
    .O(inst82_O)
  );

  //Wire declarations for instance 'inst83' (Module and_wrapped)
  wire  inst83_I0;
  wire  inst83_I1;
  wire  inst83_O;
  and_wrapped inst83(
    .I0(inst83_I0),
    .I1(inst83_I1),
    .O(inst83_O)
  );

  //Wire declarations for instance 'inst84' (Module and_wrapped)
  wire  inst84_I0;
  wire  inst84_I1;
  wire  inst84_O;
  and_wrapped inst84(
    .I0(inst84_I0),
    .I1(inst84_I1),
    .O(inst84_O)
  );

  //Wire declarations for instance 'inst85' (Module and_wrapped)
  wire  inst85_I0;
  wire  inst85_I1;
  wire  inst85_O;
  and_wrapped inst85(
    .I0(inst85_I0),
    .I1(inst85_I1),
    .O(inst85_O)
  );

  //Wire declarations for instance 'inst86' (Module and_wrapped)
  wire  inst86_I0;
  wire  inst86_I1;
  wire  inst86_O;
  and_wrapped inst86(
    .I0(inst86_I0),
    .I1(inst86_I1),
    .O(inst86_O)
  );

  //Wire declarations for instance 'inst87' (Module and_wrapped)
  wire  inst87_I0;
  wire  inst87_I1;
  wire  inst87_O;
  and_wrapped inst87(
    .I0(inst87_I0),
    .I1(inst87_I1),
    .O(inst87_O)
  );

  //Wire declarations for instance 'inst88' (Module and_wrapped)
  wire  inst88_I0;
  wire  inst88_I1;
  wire  inst88_O;
  and_wrapped inst88(
    .I0(inst88_I0),
    .I1(inst88_I1),
    .O(inst88_O)
  );

  //Wire declarations for instance 'inst89' (Module and_wrapped)
  wire  inst89_I0;
  wire  inst89_I1;
  wire  inst89_O;
  and_wrapped inst89(
    .I0(inst89_I0),
    .I1(inst89_I1),
    .O(inst89_O)
  );

  //Wire declarations for instance 'inst9' (Module and2_wrapped)
  wire [1:0] inst9_I0;
  wire [1:0] inst9_I1;
  wire [1:0] inst9_O;
  and2_wrapped inst9(
    .I0(inst9_I0),
    .I1(inst9_I1),
    .O(inst9_O)
  );

  //Wire declarations for instance 'inst90' (Module and_wrapped)
  wire  inst90_I0;
  wire  inst90_I1;
  wire  inst90_O;
  and_wrapped inst90(
    .I0(inst90_I0),
    .I1(inst90_I1),
    .O(inst90_O)
  );

  //Wire declarations for instance 'inst91' (Module fold_or8None)
  wire  inst91_I0;
  wire  inst91_I3;
  wire  inst91_O;
  wire  inst91_I4;
  wire  inst91_I2;
  wire  inst91_I1;
  wire  inst91_I7;
  wire  inst91_I5;
  wire  inst91_I6;
  fold_or8None inst91(
    .I0(inst91_I0),
    .I1(inst91_I1),
    .I2(inst91_I2),
    .I3(inst91_I3),
    .I4(inst91_I4),
    .I5(inst91_I5),
    .I6(inst91_I6),
    .I7(inst91_I7),
    .O(inst91_O)
  );

  //Wire declarations for instance 'inst92' (Module and_wrapped)
  wire  inst92_I0;
  wire  inst92_I1;
  wire  inst92_O;
  and_wrapped inst92(
    .I0(inst92_I0),
    .I1(inst92_I1),
    .O(inst92_O)
  );

  //Wire declarations for instance 'inst93' (Module and_wrapped)
  wire  inst93_I0;
  wire  inst93_I1;
  wire  inst93_O;
  and_wrapped inst93(
    .I0(inst93_I0),
    .I1(inst93_I1),
    .O(inst93_O)
  );

  //Wire declarations for instance 'inst94' (Module and_wrapped)
  wire  inst94_I0;
  wire  inst94_I1;
  wire  inst94_O;
  and_wrapped inst94(
    .I0(inst94_I0),
    .I1(inst94_I1),
    .O(inst94_O)
  );

  //Wire declarations for instance 'inst95' (Module and_wrapped)
  wire  inst95_I0;
  wire  inst95_I1;
  wire  inst95_O;
  and_wrapped inst95(
    .I0(inst95_I0),
    .I1(inst95_I1),
    .O(inst95_O)
  );

  //Wire declarations for instance 'inst96' (Module and_wrapped)
  wire  inst96_I0;
  wire  inst96_I1;
  wire  inst96_O;
  and_wrapped inst96(
    .I0(inst96_I0),
    .I1(inst96_I1),
    .O(inst96_O)
  );

  //Wire declarations for instance 'inst97' (Module and_wrapped)
  wire  inst97_I0;
  wire  inst97_I1;
  wire  inst97_O;
  and_wrapped inst97(
    .I0(inst97_I0),
    .I1(inst97_I1),
    .O(inst97_O)
  );

  //Wire declarations for instance 'inst98' (Module and_wrapped)
  wire  inst98_I0;
  wire  inst98_I1;
  wire  inst98_O;
  and_wrapped inst98(
    .I0(inst98_I0),
    .I1(inst98_I1),
    .O(inst98_O)
  );

  //Wire declarations for instance 'inst99' (Module and_wrapped)
  wire  inst99_I0;
  wire  inst99_I1;
  wire  inst99_O;
  and_wrapped inst99(
    .I0(inst99_I0),
    .I1(inst99_I1),
    .O(inst99_O)
  );

  //Wire declarations for instance 'prev_empty' (Module DFF_init1_has_ceFalse_has_resetFalse)
  wire  prev_empty_CLK;
  wire  prev_empty_I;
  wire  prev_empty_O;
  DFF_init1_has_ceFalse_has_resetFalse prev_empty(
    .CLK(prev_empty_CLK),
    .I(prev_empty_I),
    .O(prev_empty_O)
  );

  //Wire declarations for instance 'prev_full' (Module DFF_init0_has_ceFalse_has_resetFalse)
  wire  prev_full_CLK;
  wire  prev_full_I;
  wire  prev_full_O;
  DFF_init0_has_ceFalse_has_resetFalse prev_full(
    .CLK(prev_full_CLK),
    .I(prev_full_I),
    .O(prev_full_O)
  );

  //All the connections
  assign inst102_I1 = bit_const_GND_out;
  assign inst106_I1 = bit_const_GND_out;
  assign inst73_I1 = bit_const_GND_out;
  assign inst75_I1 = bit_const_GND_out;
  assign inst77_I1 = bit_const_GND_out;
  assign inst79_I1 = bit_const_GND_out;
  assign inst84_I1 = bit_const_GND_out;
  assign inst88_I1 = bit_const_GND_out;
  assign inst92_I1 = bit_const_GND_out;
  assign inst94_I1 = bit_const_GND_out;
  assign inst96_I1 = bit_const_GND_out;
  assign inst98_I1 = bit_const_GND_out;
  assign inst10_I1[0] = bit_const_GND_out;
  assign inst125_I1[1] = bit_const_GND_out;
  assign inst130_I1[1] = bit_const_GND_out;
  assign inst140_I1[1] = bit_const_GND_out;
  assign inst153_I1[1] = bit_const_GND_out;
  assign inst171_I1[1] = bit_const_GND_out;
  assign inst176_I1[1] = bit_const_GND_out;
  assign inst186_I1[1] = bit_const_GND_out;
  assign inst199_I1[1] = bit_const_GND_out;
  assign inst3_I1[0] = bit_const_GND_out;
  assign inst4_I1[0] = bit_const_GND_out;
  assign inst5_I1[0] = bit_const_GND_out;
  assign inst6_I1[0] = bit_const_GND_out;
  assign inst7_I1[0] = bit_const_GND_out;
  assign inst8_I1[0] = bit_const_GND_out;
  assign inst9_I1[0] = bit_const_GND_out;
  assign inst10_I1[1] = bit_const_VCC_out;
  assign inst125_I1[0] = bit_const_VCC_out;
  assign inst130_I1[0] = bit_const_VCC_out;
  assign inst140_I1[0] = bit_const_VCC_out;
  assign inst153_I1[0] = bit_const_VCC_out;
  assign inst171_I1[0] = bit_const_VCC_out;
  assign inst176_I1[0] = bit_const_VCC_out;
  assign inst186_I1[0] = bit_const_VCC_out;
  assign inst199_I1[0] = bit_const_VCC_out;
  assign inst3_I1[1] = bit_const_VCC_out;
  assign inst4_I1[1] = bit_const_VCC_out;
  assign inst5_I1[1] = bit_const_VCC_out;
  assign inst6_I1[1] = bit_const_VCC_out;
  assign inst7_I1[1] = bit_const_VCC_out;
  assign inst8_I1[1] = bit_const_VCC_out;
  assign inst9_I1[1] = bit_const_VCC_out;
  assign inst1_CLK = CLK;
  assign inst1_I[1:0] = inst2_O[1:0];
  assign inst2_I7[1:0] = inst10_O[1:0];
  assign inst100_I0 = inst101_O;
  assign inst100_I1 = inst102_O;
  assign inst100_I2 = inst103_O;
  assign inst100_I3 = inst104_O;
  assign inst100_I4 = inst105_O;
  assign inst100_I5 = inst106_O;
  assign inst100_I6 = inst107_O;
  assign inst100_I7 = inst108_O;
  assign empty = inst100_O;
  assign inst101_I0 = inst0_O[0];
  assign inst101_I1 = inst131_O;
  assign inst102_I0 = inst0_O[1];
  assign inst103_I0 = inst0_O[2];
  assign inst103_I1 = inst154_O;
  assign inst104_I0 = inst0_O[3];
  assign inst104_I1 = prev_empty_O;
  assign inst105_I0 = inst0_O[4];
  assign inst105_I1 = inst177_O;
  assign inst106_I0 = inst0_O[5];
  assign inst107_I0 = inst0_O[6];
  assign inst107_I1 = inst200_O;
  assign inst108_I0 = inst0_O[7];
  assign inst108_I1 = prev_empty_O;
  assign inst109_I0[3:0] = inst110_O[3:0];
  assign inst109_I1[3:0] = inst111_O[3:0];
  assign inst109_I2[3:0] = inst112_O[3:0];
  assign inst109_I3[3:0] = inst113_O[3:0];
  assign inst109_I4[3:0] = inst114_O[3:0];
  assign inst109_I5[3:0] = inst115_O[3:0];
  assign inst109_I6[3:0] = inst116_O[3:0];
  assign inst109_I7[3:0] = inst117_O[3:0];
  assign rdata[3:0] = inst109_O[3:0];
  assign inst11_CLK = CLK;
  assign inst11_I[3:0] = inst15_O[3:0];
  assign inst121_I0[3:0] = inst11_O[3:0];
  assign inst136_I0[3:0] = inst11_O[3:0];
  assign inst150_I0[3:0] = inst11_O[3:0];
  assign inst159_I0[3:0] = inst11_O[3:0];
  assign inst167_I0[3:0] = inst11_O[3:0];
  assign inst182_I0[3:0] = inst11_O[3:0];
  assign inst196_I0[3:0] = inst11_O[3:0];
  assign inst205_I0[3:0] = inst11_O[3:0];
  assign inst27_I1[3:0] = inst11_O[3:0];
  assign inst31_I1[3:0] = inst11_O[3:0];
  assign inst43_I1[3:0] = inst11_O[3:0];
  assign inst47_I1[3:0] = inst11_O[3:0];
  assign inst110_I1[3:0] = inst127_O[3:0];
  assign inst111_I1[3:0] = inst142_O[3:0];
  assign inst112_I1[3:0] = inst150_O[3:0];
  assign inst113_I1[3:0] = inst159_O[3:0];
  assign inst114_I1[3:0] = inst173_O[3:0];
  assign inst115_I1[3:0] = inst188_O[3:0];
  assign inst116_I1[3:0] = inst196_O[3:0];
  assign inst117_I1[3:0] = inst205_O[3:0];
  assign inst118_in = prev_full_O;
  assign inst119_I1 = inst118_out;
  assign inst119_I0 = wen;
  assign inst132_I1 = inst119_O;
  assign inst12_CLK = CLK;
  assign inst12_I[3:0] = inst16_O[3:0];
  assign inst122_I0[3:0] = inst12_O[3:0];
  assign inst137_I0[3:0] = inst12_O[3:0];
  assign inst150_I1[3:0] = inst12_O[3:0];
  assign inst159_I1[3:0] = inst12_O[3:0];
  assign inst168_I0[3:0] = inst12_O[3:0];
  assign inst183_I0[3:0] = inst12_O[3:0];
  assign inst196_I1[3:0] = inst12_O[3:0];
  assign inst205_I1[3:0] = inst12_O[3:0];
  assign inst28_I1[3:0] = inst12_O[3:0];
  assign inst32_I1[3:0] = inst12_O[3:0];
  assign inst44_I1[3:0] = inst12_O[3:0];
  assign inst48_I1[3:0] = inst12_O[3:0];
  assign inst120_I[1:0] = inst61_O[1:0];
  assign inst121_I1[3:0] = wdata[3:0];
  assign inst127_I0[3:0] = inst121_O[3:0];
  assign inst19_I1[3:0] = inst121_O[3:0];
  assign inst121_S = inst120_O[0];
  assign inst122_I1[3:0] = wdata[3:0];
  assign inst127_I1[3:0] = inst122_O[3:0];
  assign inst20_I1[3:0] = inst122_O[3:0];
  assign inst122_S = inst120_O[1];
  assign inst123_I0[3:0] = inst13_O[3:0];
  assign inst123_I1[3:0] = wdata[3:0];
  assign inst127_I2[3:0] = inst123_O[3:0];
  assign inst21_I1[3:0] = inst123_O[3:0];
  assign inst123_S = inst120_O[2];
  assign inst124_I0[3:0] = inst14_O[3:0];
  assign inst124_I1[3:0] = wdata[3:0];
  assign inst127_I3[3:0] = inst124_O[3:0];
  assign inst22_I1[3:0] = inst124_O[3:0];
  assign inst124_S = inst120_O[3];
  assign inst125_I0[1:0] = inst61_O[1:0];
  assign inst126_I1[1:0] = inst125_O[1:0];
  assign inst131_I1[1:0] = inst125_O[1:0];
  assign inst63_I1[1:0] = inst125_O[1:0];
  assign inst126_I0[1:0] = inst51_O[1:0];
  assign inst127_S[1:0] = inst51_O[1:0];
  assign inst128_in = prev_empty_O;
  assign inst129_I1 = inst128_out;
  assign inst129_I0 = ren;
  assign inst132_I2 = inst129_O;
  assign inst13_CLK = CLK;
  assign inst13_I[3:0] = inst17_O[3:0];
  assign inst138_I0[3:0] = inst13_O[3:0];
  assign inst150_I2[3:0] = inst13_O[3:0];
  assign inst159_I2[3:0] = inst13_O[3:0];
  assign inst169_I0[3:0] = inst13_O[3:0];
  assign inst184_I0[3:0] = inst13_O[3:0];
  assign inst196_I2[3:0] = inst13_O[3:0];
  assign inst205_I2[3:0] = inst13_O[3:0];
  assign inst29_I1[3:0] = inst13_O[3:0];
  assign inst33_I1[3:0] = inst13_O[3:0];
  assign inst45_I1[3:0] = inst13_O[3:0];
  assign inst49_I1[3:0] = inst13_O[3:0];
  assign inst130_I0[1:0] = inst51_O[1:0];
  assign inst131_I0[1:0] = inst130_O[1:0];
  assign inst53_I1[1:0] = inst130_O[1:0];
  assign inst83_I1 = inst131_O;
  assign inst132_I0 = inst1_O[0];
  assign inst0_I[0] = inst132_O;
  assign inst133_in = prev_full_O;
  assign inst134_I1 = inst133_out;
  assign inst134_I0 = wen;
  assign inst146_I1 = inst134_O;
  assign inst135_I[1:0] = inst61_O[1:0];
  assign inst136_I1[3:0] = wdata[3:0];
  assign inst142_I0[3:0] = inst136_O[3:0];
  assign inst23_I1[3:0] = inst136_O[3:0];
  assign inst136_S = inst135_O[0];
  assign inst137_I1[3:0] = wdata[3:0];
  assign inst142_I1[3:0] = inst137_O[3:0];
  assign inst24_I1[3:0] = inst137_O[3:0];
  assign inst137_S = inst135_O[1];
  assign inst138_I1[3:0] = wdata[3:0];
  assign inst142_I2[3:0] = inst138_O[3:0];
  assign inst25_I1[3:0] = inst138_O[3:0];
  assign inst138_S = inst135_O[2];
  assign inst139_I0[3:0] = inst14_O[3:0];
  assign inst139_I1[3:0] = wdata[3:0];
  assign inst142_I3[3:0] = inst139_O[3:0];
  assign inst26_I1[3:0] = inst139_O[3:0];
  assign inst139_S = inst135_O[3];
  assign inst14_CLK = CLK;
  assign inst14_I[3:0] = inst18_O[3:0];
  assign inst150_I3[3:0] = inst14_O[3:0];
  assign inst159_I3[3:0] = inst14_O[3:0];
  assign inst170_I0[3:0] = inst14_O[3:0];
  assign inst185_I0[3:0] = inst14_O[3:0];
  assign inst196_I3[3:0] = inst14_O[3:0];
  assign inst205_I3[3:0] = inst14_O[3:0];
  assign inst30_I1[3:0] = inst14_O[3:0];
  assign inst34_I1[3:0] = inst14_O[3:0];
  assign inst46_I1[3:0] = inst14_O[3:0];
  assign inst50_I1[3:0] = inst14_O[3:0];
  assign inst140_I0[1:0] = inst61_O[1:0];
  assign inst141_I1[1:0] = inst140_O[1:0];
  assign inst64_I1[1:0] = inst140_O[1:0];
  assign inst141_I0[1:0] = inst51_O[1:0];
  assign inst74_I1 = inst141_O;
  assign inst93_I1 = inst141_O;
  assign inst142_S[1:0] = inst51_O[1:0];
  assign inst143_in = prev_empty_O;
  assign inst144_I1 = inst143_out;
  assign inst144_I0 = ren;
  assign inst145_in = inst144_O;
  assign inst146_I2 = inst145_out;
  assign inst146_I0 = inst1_O[0];
  assign inst0_I[1] = inst146_O;
  assign inst147_in = prev_full_O;
  assign inst148_I1 = inst147_out;
  assign inst148_I0 = wen;
  assign inst149_in = inst148_O;
  assign inst155_I1 = inst149_out;
  assign inst15_I0[3:0] = inst19_O[3:0];
  assign inst15_I1[3:0] = inst23_O[3:0];
  assign inst15_I2[3:0] = inst27_O[3:0];
  assign inst15_I3[3:0] = inst31_O[3:0];
  assign inst15_I4[3:0] = inst35_O[3:0];
  assign inst15_I5[3:0] = inst39_O[3:0];
  assign inst15_I6[3:0] = inst43_O[3:0];
  assign inst15_I7[3:0] = inst47_O[3:0];
  assign inst150_S[1:0] = inst51_O[1:0];
  assign inst151_in = prev_empty_O;
  assign inst152_I1 = inst151_out;
  assign inst152_I0 = ren;
  assign inst155_I2 = inst152_O;
  assign inst153_I0[1:0] = inst51_O[1:0];
  assign inst154_I0[1:0] = inst153_O[1:0];
  assign inst55_I1[1:0] = inst153_O[1:0];
  assign inst154_I1[1:0] = inst61_O[1:0];
  assign inst85_I1 = inst154_O;
  assign inst155_I0 = inst1_O[0];
  assign inst0_I[2] = inst155_O;
  assign inst156_in = prev_full_O;
  assign inst157_I1 = inst156_out;
  assign inst157_I0 = wen;
  assign inst158_in = inst157_O;
  assign inst163_I1 = inst158_out;
  assign inst159_S[1:0] = inst51_O[1:0];
  assign inst16_I0[3:0] = inst20_O[3:0];
  assign inst16_I1[3:0] = inst24_O[3:0];
  assign inst16_I2[3:0] = inst28_O[3:0];
  assign inst16_I3[3:0] = inst32_O[3:0];
  assign inst16_I4[3:0] = inst36_O[3:0];
  assign inst16_I5[3:0] = inst40_O[3:0];
  assign inst16_I6[3:0] = inst44_O[3:0];
  assign inst16_I7[3:0] = inst48_O[3:0];
  assign inst160_in = prev_empty_O;
  assign inst161_I1 = inst160_out;
  assign inst161_I0 = ren;
  assign inst162_in = inst161_O;
  assign inst163_I2 = inst162_out;
  assign inst163_I0 = inst1_O[0];
  assign inst0_I[3] = inst163_O;
  assign inst164_in = prev_full_O;
  assign inst165_I1 = inst164_out;
  assign inst165_I0 = wen;
  assign inst178_I1 = inst165_O;
  assign inst166_I[1:0] = inst61_O[1:0];
  assign inst167_I1[3:0] = wdata[3:0];
  assign inst173_I0[3:0] = inst167_O[3:0];
  assign inst35_I1[3:0] = inst167_O[3:0];
  assign inst167_S = inst166_O[0];
  assign inst168_I1[3:0] = wdata[3:0];
  assign inst173_I1[3:0] = inst168_O[3:0];
  assign inst36_I1[3:0] = inst168_O[3:0];
  assign inst168_S = inst166_O[1];
  assign inst169_I1[3:0] = wdata[3:0];
  assign inst173_I2[3:0] = inst169_O[3:0];
  assign inst37_I1[3:0] = inst169_O[3:0];
  assign inst169_S = inst166_O[2];
  assign inst17_I0[3:0] = inst21_O[3:0];
  assign inst17_I1[3:0] = inst25_O[3:0];
  assign inst17_I2[3:0] = inst29_O[3:0];
  assign inst17_I3[3:0] = inst33_O[3:0];
  assign inst17_I4[3:0] = inst37_O[3:0];
  assign inst17_I5[3:0] = inst41_O[3:0];
  assign inst17_I6[3:0] = inst45_O[3:0];
  assign inst17_I7[3:0] = inst49_O[3:0];
  assign inst170_I1[3:0] = wdata[3:0];
  assign inst173_I3[3:0] = inst170_O[3:0];
  assign inst38_I1[3:0] = inst170_O[3:0];
  assign inst170_S = inst166_O[3];
  assign inst171_I0[1:0] = inst61_O[1:0];
  assign inst172_I1[1:0] = inst171_O[1:0];
  assign inst177_I1[1:0] = inst171_O[1:0];
  assign inst67_I1[1:0] = inst171_O[1:0];
  assign inst172_I0[1:0] = inst51_O[1:0];
  assign inst173_S[1:0] = inst51_O[1:0];
  assign inst174_in = prev_empty_O;
  assign inst175_I1 = inst174_out;
  assign inst175_I0 = ren;
  assign inst178_I2 = inst175_O;
  assign inst176_I0[1:0] = inst51_O[1:0];
  assign inst177_I0[1:0] = inst176_O[1:0];
  assign inst57_I1[1:0] = inst176_O[1:0];
  assign inst87_I1 = inst177_O;
  assign inst178_I0 = inst1_O[1];
  assign inst0_I[4] = inst178_O;
  assign inst179_in = prev_full_O;
  assign inst180_I1 = inst179_out;
  assign inst18_I0[3:0] = inst22_O[3:0];
  assign inst18_I1[3:0] = inst26_O[3:0];
  assign inst18_I2[3:0] = inst30_O[3:0];
  assign inst18_I3[3:0] = inst34_O[3:0];
  assign inst18_I4[3:0] = inst38_O[3:0];
  assign inst18_I5[3:0] = inst42_O[3:0];
  assign inst18_I6[3:0] = inst46_O[3:0];
  assign inst18_I7[3:0] = inst50_O[3:0];
  assign inst180_I0 = wen;
  assign inst192_I1 = inst180_O;
  assign inst181_I[1:0] = inst61_O[1:0];
  assign inst182_I1[3:0] = wdata[3:0];
  assign inst188_I0[3:0] = inst182_O[3:0];
  assign inst39_I1[3:0] = inst182_O[3:0];
  assign inst182_S = inst181_O[0];
  assign inst183_I1[3:0] = wdata[3:0];
  assign inst188_I1[3:0] = inst183_O[3:0];
  assign inst40_I1[3:0] = inst183_O[3:0];
  assign inst183_S = inst181_O[1];
  assign inst184_I1[3:0] = wdata[3:0];
  assign inst188_I2[3:0] = inst184_O[3:0];
  assign inst41_I1[3:0] = inst184_O[3:0];
  assign inst184_S = inst181_O[2];
  assign inst185_I1[3:0] = wdata[3:0];
  assign inst188_I3[3:0] = inst185_O[3:0];
  assign inst42_I1[3:0] = inst185_O[3:0];
  assign inst185_S = inst181_O[3];
  assign inst186_I0[1:0] = inst61_O[1:0];
  assign inst187_I1[1:0] = inst186_O[1:0];
  assign inst68_I1[1:0] = inst186_O[1:0];
  assign inst187_I0[1:0] = inst51_O[1:0];
  assign inst78_I1 = inst187_O;
  assign inst97_I1 = inst187_O;
  assign inst188_S[1:0] = inst51_O[1:0];
  assign inst189_in = prev_empty_O;
  assign inst190_I1 = inst189_out;
  assign inst190_I0 = ren;
  assign inst191_in = inst190_O;
  assign inst192_I2 = inst191_out;
  assign inst192_I0 = inst1_O[1];
  assign inst0_I[5] = inst192_O;
  assign inst193_in = prev_full_O;
  assign inst194_I1 = inst193_out;
  assign inst194_I0 = wen;
  assign inst195_in = inst194_O;
  assign inst201_I1 = inst195_out;
  assign inst196_S[1:0] = inst51_O[1:0];
  assign inst197_in = prev_empty_O;
  assign inst198_I1 = inst197_out;
  assign inst198_I0 = ren;
  assign inst201_I2 = inst198_O;
  assign inst199_I0[1:0] = inst51_O[1:0];
  assign inst200_I0[1:0] = inst199_O[1:0];
  assign inst59_I1[1:0] = inst199_O[1:0];
  assign inst2_I0[1:0] = inst3_O[1:0];
  assign inst2_I1[1:0] = inst4_O[1:0];
  assign inst2_I2[1:0] = inst5_O[1:0];
  assign inst2_I3[1:0] = inst6_O[1:0];
  assign inst2_I4[1:0] = inst7_O[1:0];
  assign inst2_I5[1:0] = inst8_O[1:0];
  assign inst2_I6[1:0] = inst9_O[1:0];
  assign inst200_I1[1:0] = inst61_O[1:0];
  assign inst89_I1 = inst200_O;
  assign inst201_I0 = inst1_O[1];
  assign inst0_I[6] = inst201_O;
  assign inst202_in = prev_full_O;
  assign inst203_I1 = inst202_out;
  assign inst203_I0 = wen;
  assign inst204_in = inst203_O;
  assign inst209_I1 = inst204_out;
  assign inst205_S[1:0] = inst51_O[1:0];
  assign inst206_in = prev_empty_O;
  assign inst207_I1 = inst206_out;
  assign inst207_I0 = ren;
  assign inst208_in = inst207_O;
  assign inst209_I2 = inst208_out;
  assign inst209_I0 = inst1_O[1];
  assign inst0_I[7] = inst209_O;
  assign inst51_CLK = CLK;
  assign inst51_I[1:0] = inst52_O[1:0];
  assign inst54_I1[1:0] = inst51_O[1:0];
  assign inst56_I1[1:0] = inst51_O[1:0];
  assign inst58_I1[1:0] = inst51_O[1:0];
  assign inst60_I1[1:0] = inst51_O[1:0];
  assign inst52_I0[1:0] = inst53_O[1:0];
  assign inst52_I1[1:0] = inst54_O[1:0];
  assign inst52_I2[1:0] = inst55_O[1:0];
  assign inst52_I3[1:0] = inst56_O[1:0];
  assign inst52_I4[1:0] = inst57_O[1:0];
  assign inst52_I5[1:0] = inst58_O[1:0];
  assign inst52_I6[1:0] = inst59_O[1:0];
  assign inst52_I7[1:0] = inst60_O[1:0];
  assign inst61_CLK = CLK;
  assign inst61_I[1:0] = inst62_O[1:0];
  assign inst65_I1[1:0] = inst61_O[1:0];
  assign inst66_I1[1:0] = inst61_O[1:0];
  assign inst69_I1[1:0] = inst61_O[1:0];
  assign inst70_I1[1:0] = inst61_O[1:0];
  assign inst62_I0[1:0] = inst63_O[1:0];
  assign inst62_I1[1:0] = inst64_O[1:0];
  assign inst62_I2[1:0] = inst65_O[1:0];
  assign inst62_I3[1:0] = inst66_O[1:0];
  assign inst62_I4[1:0] = inst67_O[1:0];
  assign inst62_I5[1:0] = inst68_O[1:0];
  assign inst62_I6[1:0] = inst69_O[1:0];
  assign inst62_I7[1:0] = inst70_O[1:0];
  assign inst72_I0 = inst73_O;
  assign inst72_I1 = inst74_O;
  assign inst72_I2 = inst75_O;
  assign inst72_I3 = inst76_O;
  assign inst72_I4 = inst77_O;
  assign inst72_I5 = inst78_O;
  assign inst72_I6 = inst79_O;
  assign inst72_I7 = inst80_O;
  assign prev_full_I = inst72_O;
  assign inst73_I0 = inst0_O[0];
  assign inst74_I0 = inst0_O[1];
  assign inst75_I0 = inst0_O[2];
  assign inst76_I0 = inst0_O[3];
  assign inst76_I1 = prev_full_O;
  assign inst77_I0 = inst0_O[4];
  assign inst78_I0 = inst0_O[5];
  assign inst79_I0 = inst0_O[6];
  assign inst80_I0 = inst0_O[7];
  assign inst80_I1 = prev_full_O;
  assign inst82_I0 = inst83_O;
  assign inst82_I1 = inst84_O;
  assign inst82_I2 = inst85_O;
  assign inst82_I3 = inst86_O;
  assign inst82_I4 = inst87_O;
  assign inst82_I5 = inst88_O;
  assign inst82_I6 = inst89_O;
  assign inst82_I7 = inst90_O;
  assign prev_empty_I = inst82_O;
  assign inst83_I0 = inst0_O[0];
  assign inst84_I0 = inst0_O[1];
  assign inst85_I0 = inst0_O[2];
  assign inst86_I0 = inst0_O[3];
  assign inst86_I1 = prev_empty_O;
  assign inst87_I0 = inst0_O[4];
  assign inst88_I0 = inst0_O[5];
  assign inst89_I0 = inst0_O[6];
  assign inst90_I0 = inst0_O[7];
  assign inst90_I1 = prev_empty_O;
  assign inst91_I0 = inst92_O;
  assign inst91_I1 = inst93_O;
  assign inst91_I2 = inst94_O;
  assign inst91_I3 = inst95_O;
  assign inst91_I4 = inst96_O;
  assign inst91_I5 = inst97_O;
  assign inst91_I6 = inst98_O;
  assign inst91_I7 = inst99_O;
  assign full = inst91_O;
  assign inst92_I0 = inst0_O[0];
  assign inst93_I0 = inst0_O[1];
  assign inst94_I0 = inst0_O[2];
  assign inst95_I0 = inst0_O[3];
  assign inst95_I1 = prev_full_O;
  assign inst96_I0 = inst0_O[4];
  assign inst97_I0 = inst0_O[5];
  assign inst98_I0 = inst0_O[6];
  assign inst99_I0 = inst0_O[7];
  assign inst99_I1 = prev_full_O;
  assign prev_empty_CLK = CLK;
  assign prev_full_CLK = CLK;
  assign inst110_I0[0] = inst0_O[0];
  assign inst110_I0[1] = inst0_O[0];
  assign inst110_I0[2] = inst0_O[0];
  assign inst110_I0[3] = inst0_O[0];
  assign inst19_I0[0] = inst0_O[0];
  assign inst19_I0[1] = inst0_O[0];
  assign inst19_I0[2] = inst0_O[0];
  assign inst19_I0[3] = inst0_O[0];
  assign inst20_I0[0] = inst0_O[0];
  assign inst20_I0[1] = inst0_O[0];
  assign inst20_I0[2] = inst0_O[0];
  assign inst20_I0[3] = inst0_O[0];
  assign inst21_I0[0] = inst0_O[0];
  assign inst21_I0[1] = inst0_O[0];
  assign inst21_I0[2] = inst0_O[0];
  assign inst21_I0[3] = inst0_O[0];
  assign inst22_I0[0] = inst0_O[0];
  assign inst22_I0[1] = inst0_O[0];
  assign inst22_I0[2] = inst0_O[0];
  assign inst22_I0[3] = inst0_O[0];
  assign inst3_I0[0] = inst0_O[0];
  assign inst3_I0[1] = inst0_O[0];
  assign inst53_I0[0] = inst0_O[0];
  assign inst53_I0[1] = inst0_O[0];
  assign inst63_I0[0] = inst0_O[0];
  assign inst63_I0[1] = inst0_O[0];
  assign inst111_I0[0] = inst0_O[1];
  assign inst111_I0[1] = inst0_O[1];
  assign inst111_I0[2] = inst0_O[1];
  assign inst111_I0[3] = inst0_O[1];
  assign inst23_I0[0] = inst0_O[1];
  assign inst23_I0[1] = inst0_O[1];
  assign inst23_I0[2] = inst0_O[1];
  assign inst23_I0[3] = inst0_O[1];
  assign inst24_I0[0] = inst0_O[1];
  assign inst24_I0[1] = inst0_O[1];
  assign inst24_I0[2] = inst0_O[1];
  assign inst24_I0[3] = inst0_O[1];
  assign inst25_I0[0] = inst0_O[1];
  assign inst25_I0[1] = inst0_O[1];
  assign inst25_I0[2] = inst0_O[1];
  assign inst25_I0[3] = inst0_O[1];
  assign inst26_I0[0] = inst0_O[1];
  assign inst26_I0[1] = inst0_O[1];
  assign inst26_I0[2] = inst0_O[1];
  assign inst26_I0[3] = inst0_O[1];
  assign inst4_I0[0] = inst0_O[1];
  assign inst4_I0[1] = inst0_O[1];
  assign inst54_I0[0] = inst0_O[1];
  assign inst54_I0[1] = inst0_O[1];
  assign inst64_I0[0] = inst0_O[1];
  assign inst64_I0[1] = inst0_O[1];
  assign inst112_I0[0] = inst0_O[2];
  assign inst112_I0[1] = inst0_O[2];
  assign inst112_I0[2] = inst0_O[2];
  assign inst112_I0[3] = inst0_O[2];
  assign inst27_I0[0] = inst0_O[2];
  assign inst27_I0[1] = inst0_O[2];
  assign inst27_I0[2] = inst0_O[2];
  assign inst27_I0[3] = inst0_O[2];
  assign inst28_I0[0] = inst0_O[2];
  assign inst28_I0[1] = inst0_O[2];
  assign inst28_I0[2] = inst0_O[2];
  assign inst28_I0[3] = inst0_O[2];
  assign inst29_I0[0] = inst0_O[2];
  assign inst29_I0[1] = inst0_O[2];
  assign inst29_I0[2] = inst0_O[2];
  assign inst29_I0[3] = inst0_O[2];
  assign inst30_I0[0] = inst0_O[2];
  assign inst30_I0[1] = inst0_O[2];
  assign inst30_I0[2] = inst0_O[2];
  assign inst30_I0[3] = inst0_O[2];
  assign inst5_I0[0] = inst0_O[2];
  assign inst5_I0[1] = inst0_O[2];
  assign inst55_I0[0] = inst0_O[2];
  assign inst55_I0[1] = inst0_O[2];
  assign inst65_I0[0] = inst0_O[2];
  assign inst65_I0[1] = inst0_O[2];
  assign inst113_I0[0] = inst0_O[3];
  assign inst113_I0[1] = inst0_O[3];
  assign inst113_I0[2] = inst0_O[3];
  assign inst113_I0[3] = inst0_O[3];
  assign inst31_I0[0] = inst0_O[3];
  assign inst31_I0[1] = inst0_O[3];
  assign inst31_I0[2] = inst0_O[3];
  assign inst31_I0[3] = inst0_O[3];
  assign inst32_I0[0] = inst0_O[3];
  assign inst32_I0[1] = inst0_O[3];
  assign inst32_I0[2] = inst0_O[3];
  assign inst32_I0[3] = inst0_O[3];
  assign inst33_I0[0] = inst0_O[3];
  assign inst33_I0[1] = inst0_O[3];
  assign inst33_I0[2] = inst0_O[3];
  assign inst33_I0[3] = inst0_O[3];
  assign inst34_I0[0] = inst0_O[3];
  assign inst34_I0[1] = inst0_O[3];
  assign inst34_I0[2] = inst0_O[3];
  assign inst34_I0[3] = inst0_O[3];
  assign inst56_I0[0] = inst0_O[3];
  assign inst56_I0[1] = inst0_O[3];
  assign inst6_I0[0] = inst0_O[3];
  assign inst6_I0[1] = inst0_O[3];
  assign inst66_I0[0] = inst0_O[3];
  assign inst66_I0[1] = inst0_O[3];
  assign inst114_I0[0] = inst0_O[4];
  assign inst114_I0[1] = inst0_O[4];
  assign inst114_I0[2] = inst0_O[4];
  assign inst114_I0[3] = inst0_O[4];
  assign inst35_I0[0] = inst0_O[4];
  assign inst35_I0[1] = inst0_O[4];
  assign inst35_I0[2] = inst0_O[4];
  assign inst35_I0[3] = inst0_O[4];
  assign inst36_I0[0] = inst0_O[4];
  assign inst36_I0[1] = inst0_O[4];
  assign inst36_I0[2] = inst0_O[4];
  assign inst36_I0[3] = inst0_O[4];
  assign inst37_I0[0] = inst0_O[4];
  assign inst37_I0[1] = inst0_O[4];
  assign inst37_I0[2] = inst0_O[4];
  assign inst37_I0[3] = inst0_O[4];
  assign inst38_I0[0] = inst0_O[4];
  assign inst38_I0[1] = inst0_O[4];
  assign inst38_I0[2] = inst0_O[4];
  assign inst38_I0[3] = inst0_O[4];
  assign inst57_I0[0] = inst0_O[4];
  assign inst57_I0[1] = inst0_O[4];
  assign inst67_I0[0] = inst0_O[4];
  assign inst67_I0[1] = inst0_O[4];
  assign inst7_I0[0] = inst0_O[4];
  assign inst7_I0[1] = inst0_O[4];
  assign inst115_I0[0] = inst0_O[5];
  assign inst115_I0[1] = inst0_O[5];
  assign inst115_I0[2] = inst0_O[5];
  assign inst115_I0[3] = inst0_O[5];
  assign inst39_I0[0] = inst0_O[5];
  assign inst39_I0[1] = inst0_O[5];
  assign inst39_I0[2] = inst0_O[5];
  assign inst39_I0[3] = inst0_O[5];
  assign inst40_I0[0] = inst0_O[5];
  assign inst40_I0[1] = inst0_O[5];
  assign inst40_I0[2] = inst0_O[5];
  assign inst40_I0[3] = inst0_O[5];
  assign inst41_I0[0] = inst0_O[5];
  assign inst41_I0[1] = inst0_O[5];
  assign inst41_I0[2] = inst0_O[5];
  assign inst41_I0[3] = inst0_O[5];
  assign inst42_I0[0] = inst0_O[5];
  assign inst42_I0[1] = inst0_O[5];
  assign inst42_I0[2] = inst0_O[5];
  assign inst42_I0[3] = inst0_O[5];
  assign inst58_I0[0] = inst0_O[5];
  assign inst58_I0[1] = inst0_O[5];
  assign inst68_I0[0] = inst0_O[5];
  assign inst68_I0[1] = inst0_O[5];
  assign inst8_I0[0] = inst0_O[5];
  assign inst8_I0[1] = inst0_O[5];
  assign inst116_I0[0] = inst0_O[6];
  assign inst116_I0[1] = inst0_O[6];
  assign inst116_I0[2] = inst0_O[6];
  assign inst116_I0[3] = inst0_O[6];
  assign inst43_I0[0] = inst0_O[6];
  assign inst43_I0[1] = inst0_O[6];
  assign inst43_I0[2] = inst0_O[6];
  assign inst43_I0[3] = inst0_O[6];
  assign inst44_I0[0] = inst0_O[6];
  assign inst44_I0[1] = inst0_O[6];
  assign inst44_I0[2] = inst0_O[6];
  assign inst44_I0[3] = inst0_O[6];
  assign inst45_I0[0] = inst0_O[6];
  assign inst45_I0[1] = inst0_O[6];
  assign inst45_I0[2] = inst0_O[6];
  assign inst45_I0[3] = inst0_O[6];
  assign inst46_I0[0] = inst0_O[6];
  assign inst46_I0[1] = inst0_O[6];
  assign inst46_I0[2] = inst0_O[6];
  assign inst46_I0[3] = inst0_O[6];
  assign inst59_I0[0] = inst0_O[6];
  assign inst59_I0[1] = inst0_O[6];
  assign inst69_I0[0] = inst0_O[6];
  assign inst69_I0[1] = inst0_O[6];
  assign inst9_I0[0] = inst0_O[6];
  assign inst9_I0[1] = inst0_O[6];
  assign inst10_I0[0] = inst0_O[7];
  assign inst10_I0[1] = inst0_O[7];
  assign inst117_I0[0] = inst0_O[7];
  assign inst117_I0[1] = inst0_O[7];
  assign inst117_I0[2] = inst0_O[7];
  assign inst117_I0[3] = inst0_O[7];
  assign inst47_I0[0] = inst0_O[7];
  assign inst47_I0[1] = inst0_O[7];
  assign inst47_I0[2] = inst0_O[7];
  assign inst47_I0[3] = inst0_O[7];
  assign inst48_I0[0] = inst0_O[7];
  assign inst48_I0[1] = inst0_O[7];
  assign inst48_I0[2] = inst0_O[7];
  assign inst48_I0[3] = inst0_O[7];
  assign inst49_I0[0] = inst0_O[7];
  assign inst49_I0[1] = inst0_O[7];
  assign inst49_I0[2] = inst0_O[7];
  assign inst49_I0[3] = inst0_O[7];
  assign inst50_I0[0] = inst0_O[7];
  assign inst50_I0[1] = inst0_O[7];
  assign inst50_I0[2] = inst0_O[7];
  assign inst50_I0[3] = inst0_O[7];
  assign inst60_I0[0] = inst0_O[7];
  assign inst60_I0[1] = inst0_O[7];
  assign inst70_I0[0] = inst0_O[7];
  assign inst70_I0[1] = inst0_O[7];

endmodule //Fifo
