module DownsampleChannel_tb;
    wire [15:0] data_out_data;

    wire data_out_valid;

    wire data_in_ready;

    reg [15:0] data_in_data;

    reg data_in_valid;

    reg data_out_ready;

    reg CLK;


    DownsampleChannel #(
        
    ) dut (
        .data_out_data(data_out_data),
        .data_out_valid(data_out_valid),
        .data_in_ready(data_in_ready),
        .data_in_data(data_in_data),
        .data_in_valid(data_in_valid),
        .data_out_ready(data_out_ready),
        .CLK(CLK)
    );

    initial begin
        CLK = 1'd1;
        #5;
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd0;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd0)) begin
            $error("Failed on action=5 checking port data_out_data. Expected %x, got %x" , 16'd0, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd2;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd2)) begin
            $error("Failed on action=28 checking port data_out_data. Expected %x, got %x" , 16'd2, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=29 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=30 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=35 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd3;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=40 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=41 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=46 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd4;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd4)) begin
            $error("Failed on action=51 checking port data_out_data. Expected %x, got %x" , 16'd4, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=52 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=53 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=58 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd5;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=63 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=64 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=69 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd6;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd6)) begin
            $error("Failed on action=74 checking port data_out_data. Expected %x, got %x" , 16'd6, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=75 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=76 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=81 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd7;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=86 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=87 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=92 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd8;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd8)) begin
            $error("Failed on action=97 checking port data_out_data. Expected %x, got %x" , 16'd8, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=98 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=99 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd9;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=109 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=110 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd10;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd10)) begin
            $error("Failed on action=120 checking port data_out_data. Expected %x, got %x" , 16'd10, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=121 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=122 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd11;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=133 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd12;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd12)) begin
            $error("Failed on action=143 checking port data_out_data. Expected %x, got %x" , 16'd12, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=144 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=145 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd13;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=156 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=161 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd14;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd14)) begin
            $error("Failed on action=166 checking port data_out_data. Expected %x, got %x" , 16'd14, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=167 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=168 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd15;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=178 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=179 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=184 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd16;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd16)) begin
            $error("Failed on action=189 checking port data_out_data. Expected %x, got %x" , 16'd16, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=190 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=191 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd17;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=201 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=202 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=207 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd18;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd18)) begin
            $error("Failed on action=212 checking port data_out_data. Expected %x, got %x" , 16'd18, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=213 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=214 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd19;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=224 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=225 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=230 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd20;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd20)) begin
            $error("Failed on action=235 checking port data_out_data. Expected %x, got %x" , 16'd20, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=236 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=237 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd21;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=248 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd22;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd22)) begin
            $error("Failed on action=258 checking port data_out_data. Expected %x, got %x" , 16'd22, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=259 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=260 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=265 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd23;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=271 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd24;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd24)) begin
            $error("Failed on action=281 checking port data_out_data. Expected %x, got %x" , 16'd24, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=282 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=283 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=288 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd25;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=293 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=294 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=299 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd26;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd26)) begin
            $error("Failed on action=304 checking port data_out_data. Expected %x, got %x" , 16'd26, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=305 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=306 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=311 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd27;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=316 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=317 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=322 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd28;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd28)) begin
            $error("Failed on action=327 checking port data_out_data. Expected %x, got %x" , 16'd28, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=328 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=329 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=334 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd29;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=339 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=340 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=345 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd30;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd30)) begin
            $error("Failed on action=350 checking port data_out_data. Expected %x, got %x" , 16'd30, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=351 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=352 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=357 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd31;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=362 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=363 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=368 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd32;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=373 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=374 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd33;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=385 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd34;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=395 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=396 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd35;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=406 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=407 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd36;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=417 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=418 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=423 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd37;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=428 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=429 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=434 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd38;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=439 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=440 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=445 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd39;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=450 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=451 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=456 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd40;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=461 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=462 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=467 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd41;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=472 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=473 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=478 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd42;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=483 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=484 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=489 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd43;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=494 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=495 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=500 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd44;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=505 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=506 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=511 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd45;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=517 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=522 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd46;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=528 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd47;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=538 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=539 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd48;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=549 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=550 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd49;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=560 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=561 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=566 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd50;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=571 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=572 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=577 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd51;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=582 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=583 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=588 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd52;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=593 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=594 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=599 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd53;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=604 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=605 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=610 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd54;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=615 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=616 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=621 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd55;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=626 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=627 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=632 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd56;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=637 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=638 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=643 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd57;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=648 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=649 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=654 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd58;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=660 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd59;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=671 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd60;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=682 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd61;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=693 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd62;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=703 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=704 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd63;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=714 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=715 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=720 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd64;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd64)) begin
            $error("Failed on action=725 checking port data_out_data. Expected %x, got %x" , 16'd64, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=726 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=727 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd65;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=737 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=738 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=743 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd66;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd66)) begin
            $error("Failed on action=748 checking port data_out_data. Expected %x, got %x" , 16'd66, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=749 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=750 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd67;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=760 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=761 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=766 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd68;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd68)) begin
            $error("Failed on action=771 checking port data_out_data. Expected %x, got %x" , 16'd68, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=772 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=773 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd69;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=783 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=784 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=789 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd70;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd70)) begin
            $error("Failed on action=794 checking port data_out_data. Expected %x, got %x" , 16'd70, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=795 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=796 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd71;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=806 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=807 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=812 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd72;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd72)) begin
            $error("Failed on action=817 checking port data_out_data. Expected %x, got %x" , 16'd72, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=818 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=819 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd73;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=829 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=830 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd74;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd74)) begin
            $error("Failed on action=840 checking port data_out_data. Expected %x, got %x" , 16'd74, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=841 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=842 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd75;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=853 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd76;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd76)) begin
            $error("Failed on action=863 checking port data_out_data. Expected %x, got %x" , 16'd76, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=864 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=865 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd77;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=876 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=881 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd78;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd78)) begin
            $error("Failed on action=886 checking port data_out_data. Expected %x, got %x" , 16'd78, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=887 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=888 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd79;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=898 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=899 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=904 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd80;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd80)) begin
            $error("Failed on action=909 checking port data_out_data. Expected %x, got %x" , 16'd80, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=910 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=911 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd81;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=921 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=922 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=927 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd82;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd82)) begin
            $error("Failed on action=932 checking port data_out_data. Expected %x, got %x" , 16'd82, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=933 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=934 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd83;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=944 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=945 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=950 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd84;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd84)) begin
            $error("Failed on action=955 checking port data_out_data. Expected %x, got %x" , 16'd84, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=956 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=957 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd85;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=968 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd86;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd86)) begin
            $error("Failed on action=978 checking port data_out_data. Expected %x, got %x" , 16'd86, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=979 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=980 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=985 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd87;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=991 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd88;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd88)) begin
            $error("Failed on action=1001 checking port data_out_data. Expected %x, got %x" , 16'd88, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1002 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1003 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1008 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd89;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1013 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1014 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1019 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd90;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd90)) begin
            $error("Failed on action=1024 checking port data_out_data. Expected %x, got %x" , 16'd90, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1025 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1026 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1031 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd91;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1036 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1037 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1042 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd92;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd92)) begin
            $error("Failed on action=1047 checking port data_out_data. Expected %x, got %x" , 16'd92, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1048 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1049 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1054 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd93;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1059 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1060 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1065 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd94;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd94)) begin
            $error("Failed on action=1070 checking port data_out_data. Expected %x, got %x" , 16'd94, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1071 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1072 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1077 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd95;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1082 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1083 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1088 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd96;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1093 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1094 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd97;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1105 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd98;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1116 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd99;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1126 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1127 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd100;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1137 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1138 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1143 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd101;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1148 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1149 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1154 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd102;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1159 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1160 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1165 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd103;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1170 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1171 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1176 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd104;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1181 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1182 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1187 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd105;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1192 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1193 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1198 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd106;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1203 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1204 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1209 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd107;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1214 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1215 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1220 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd108;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1225 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1226 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1231 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd109;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1236 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1237 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd110;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1248 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd111;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1258 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1259 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd112;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1269 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1270 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd113;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1280 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1281 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1286 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd114;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1291 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1292 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1297 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd115;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1302 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1303 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1308 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd116;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1313 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1314 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1319 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd117;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1324 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1325 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1330 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd118;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1335 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1336 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1341 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd119;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1346 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1347 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1352 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd120;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1357 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1358 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1363 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd121;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1368 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1369 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1374 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd122;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1380 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1385 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd123;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1391 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd124;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1402 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd125;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1413 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd126;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1423 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1424 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd127;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1434 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1435 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1440 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd128;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd128)) begin
            $error("Failed on action=1445 checking port data_out_data. Expected %x, got %x" , 16'd128, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1446 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1447 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd129;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1457 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1458 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1463 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd130;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd130)) begin
            $error("Failed on action=1468 checking port data_out_data. Expected %x, got %x" , 16'd130, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1469 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1470 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd131;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1480 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1481 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1486 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd132;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd132)) begin
            $error("Failed on action=1491 checking port data_out_data. Expected %x, got %x" , 16'd132, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1492 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1493 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd133;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1503 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1504 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1509 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd134;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd134)) begin
            $error("Failed on action=1514 checking port data_out_data. Expected %x, got %x" , 16'd134, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1515 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1516 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd135;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1526 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1527 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1532 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd136;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd136)) begin
            $error("Failed on action=1537 checking port data_out_data. Expected %x, got %x" , 16'd136, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1538 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1539 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd137;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1549 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1550 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd138;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd138)) begin
            $error("Failed on action=1560 checking port data_out_data. Expected %x, got %x" , 16'd138, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1561 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1562 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd139;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1573 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd140;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd140)) begin
            $error("Failed on action=1583 checking port data_out_data. Expected %x, got %x" , 16'd140, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1584 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1585 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd141;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1595 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1596 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1601 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd142;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd142)) begin
            $error("Failed on action=1606 checking port data_out_data. Expected %x, got %x" , 16'd142, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1607 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1608 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd143;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1618 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1619 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1624 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd144;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd144)) begin
            $error("Failed on action=1629 checking port data_out_data. Expected %x, got %x" , 16'd144, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1630 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1631 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd145;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1641 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1642 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1647 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd146;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd146)) begin
            $error("Failed on action=1652 checking port data_out_data. Expected %x, got %x" , 16'd146, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1653 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1654 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd147;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1664 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1665 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd148;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd148)) begin
            $error("Failed on action=1675 checking port data_out_data. Expected %x, got %x" , 16'd148, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1676 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1677 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd149;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1688 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd150;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd150)) begin
            $error("Failed on action=1698 checking port data_out_data. Expected %x, got %x" , 16'd150, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1699 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1700 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1705 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd151;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1711 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1716 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd152;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd152)) begin
            $error("Failed on action=1721 checking port data_out_data. Expected %x, got %x" , 16'd152, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1722 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1723 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1728 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd153;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1733 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1734 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1739 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd154;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd154)) begin
            $error("Failed on action=1744 checking port data_out_data. Expected %x, got %x" , 16'd154, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1745 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1746 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1751 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd155;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1756 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1757 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1762 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd156;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd156)) begin
            $error("Failed on action=1767 checking port data_out_data. Expected %x, got %x" , 16'd156, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1768 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1769 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1774 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd157;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1779 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1780 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1785 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd158;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd158)) begin
            $error("Failed on action=1790 checking port data_out_data. Expected %x, got %x" , 16'd158, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=1791 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1792 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1797 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd159;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1802 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1803 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1808 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd160;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1813 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1814 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd161;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1825 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd162;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1836 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd163;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1846 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1847 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd164;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1857 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1858 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1863 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd165;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1868 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1869 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1874 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd166;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1879 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1880 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1885 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd167;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1890 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1891 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1896 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd168;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1901 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1902 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1907 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd169;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1912 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1913 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1918 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd170;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1923 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1924 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1929 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd171;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1934 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1935 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1940 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd172;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1945 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1946 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1951 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd173;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1956 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1957 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd174;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1968 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd175;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1978 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1979 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd176;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1989 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=1990 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=1995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd177;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2000 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2001 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2006 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd178;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2011 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2012 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2017 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd179;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2022 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2023 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2028 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd180;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2033 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2034 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2039 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd181;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2044 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2045 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2050 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd182;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2055 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2056 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2061 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd183;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2066 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2067 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2072 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd184;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2077 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2078 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2083 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd185;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2088 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2089 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2094 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd186;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2100 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2105 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd187;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2111 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd188;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2122 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd189;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2133 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd190;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2143 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2144 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2149 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd191;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2154 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2155 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2160 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd192;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd192)) begin
            $error("Failed on action=2165 checking port data_out_data. Expected %x, got %x" , 16'd192, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2166 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2167 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2172 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd193;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2177 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2178 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2183 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd194;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd194)) begin
            $error("Failed on action=2188 checking port data_out_data. Expected %x, got %x" , 16'd194, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2189 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2190 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2195 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd195;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2200 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2201 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2206 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd196;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd196)) begin
            $error("Failed on action=2211 checking port data_out_data. Expected %x, got %x" , 16'd196, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2212 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2213 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2218 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd197;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2223 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2224 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2229 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd198;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd198)) begin
            $error("Failed on action=2234 checking port data_out_data. Expected %x, got %x" , 16'd198, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2235 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2236 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2241 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd199;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2246 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2247 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2252 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd200;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd200)) begin
            $error("Failed on action=2257 checking port data_out_data. Expected %x, got %x" , 16'd200, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2258 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2259 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd201;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2269 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2270 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd202;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd202)) begin
            $error("Failed on action=2280 checking port data_out_data. Expected %x, got %x" , 16'd202, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2281 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2282 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd203;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2293 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd204;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd204)) begin
            $error("Failed on action=2303 checking port data_out_data. Expected %x, got %x" , 16'd204, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2304 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2305 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2310 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd205;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2315 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2316 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2321 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd206;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd206)) begin
            $error("Failed on action=2326 checking port data_out_data. Expected %x, got %x" , 16'd206, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2327 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2328 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2333 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd207;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2338 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2339 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2344 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd208;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd208)) begin
            $error("Failed on action=2349 checking port data_out_data. Expected %x, got %x" , 16'd208, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2350 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2351 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2356 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd209;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2361 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2362 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2367 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd210;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd210)) begin
            $error("Failed on action=2372 checking port data_out_data. Expected %x, got %x" , 16'd210, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2373 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2374 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd211;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2385 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd212;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd212)) begin
            $error("Failed on action=2395 checking port data_out_data. Expected %x, got %x" , 16'd212, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2396 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2397 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2402 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd213;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2408 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd214;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd214)) begin
            $error("Failed on action=2418 checking port data_out_data. Expected %x, got %x" , 16'd214, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2419 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2420 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2425 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd215;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2430 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2431 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2436 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd216;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd216)) begin
            $error("Failed on action=2441 checking port data_out_data. Expected %x, got %x" , 16'd216, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2442 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2443 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2448 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd217;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2453 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2454 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2459 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd218;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd218)) begin
            $error("Failed on action=2464 checking port data_out_data. Expected %x, got %x" , 16'd218, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2465 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2466 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2471 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd219;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2476 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2477 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2482 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd220;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd220)) begin
            $error("Failed on action=2487 checking port data_out_data. Expected %x, got %x" , 16'd220, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2488 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2489 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2494 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd221;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2499 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2500 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2505 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd222;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd222)) begin
            $error("Failed on action=2510 checking port data_out_data. Expected %x, got %x" , 16'd222, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2511 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2512 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2517 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd223;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2522 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2523 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2528 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd224;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2534 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd225;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2545 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd226;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2556 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd227;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2566 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2567 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd228;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2577 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2578 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2583 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd229;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2588 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2589 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2594 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd230;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2599 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2600 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2605 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd231;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2610 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2611 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2616 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd232;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2621 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2622 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2627 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd233;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2632 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2633 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2638 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd234;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2643 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2644 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2649 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd235;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2654 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2655 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2660 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd236;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2666 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2671 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd237;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2677 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd238;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2688 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd239;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2699 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd240;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2710 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd241;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2720 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2721 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2726 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd242;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2731 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2732 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2737 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd243;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2742 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2743 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2748 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd244;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2753 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2754 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2759 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd245;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2764 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2765 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2770 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd246;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2775 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2776 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2781 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd247;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2786 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2787 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2792 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd248;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2797 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2798 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2803 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd249;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2808 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2809 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2814 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd250;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2820 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2825 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd251;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2831 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd252;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2842 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd253;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2853 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd254;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2863 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2864 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2869 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd255;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2874 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2875 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2880 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd256;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd256)) begin
            $error("Failed on action=2885 checking port data_out_data. Expected %x, got %x" , 16'd256, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2886 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2887 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2892 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd257;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2897 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2898 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2903 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd258;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd258)) begin
            $error("Failed on action=2908 checking port data_out_data. Expected %x, got %x" , 16'd258, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2909 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2910 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2915 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd259;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2920 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2921 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2926 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd260;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd260)) begin
            $error("Failed on action=2931 checking port data_out_data. Expected %x, got %x" , 16'd260, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2932 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2933 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2938 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd261;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2943 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2944 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2949 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd262;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd262)) begin
            $error("Failed on action=2954 checking port data_out_data. Expected %x, got %x" , 16'd262, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2955 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2956 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2961 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd263;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2966 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2967 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2972 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd264;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd264)) begin
            $error("Failed on action=2977 checking port data_out_data. Expected %x, got %x" , 16'd264, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=2978 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2979 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd265;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2989 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=2990 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=2995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd266;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd266)) begin
            $error("Failed on action=3000 checking port data_out_data. Expected %x, got %x" , 16'd266, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3001 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3002 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd267;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3013 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd268;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd268)) begin
            $error("Failed on action=3023 checking port data_out_data. Expected %x, got %x" , 16'd268, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3024 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3025 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3030 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd269;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3035 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3036 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3041 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd270;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd270)) begin
            $error("Failed on action=3046 checking port data_out_data. Expected %x, got %x" , 16'd270, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3047 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3048 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3053 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd271;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3058 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3059 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3064 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd272;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd272)) begin
            $error("Failed on action=3069 checking port data_out_data. Expected %x, got %x" , 16'd272, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3070 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3071 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3076 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd273;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3081 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3082 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3087 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd274;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd274)) begin
            $error("Failed on action=3092 checking port data_out_data. Expected %x, got %x" , 16'd274, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3093 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3094 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd275;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3105 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd276;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd276)) begin
            $error("Failed on action=3115 checking port data_out_data. Expected %x, got %x" , 16'd276, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3116 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3117 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3122 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd277;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3128 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd278;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd278)) begin
            $error("Failed on action=3138 checking port data_out_data. Expected %x, got %x" , 16'd278, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3139 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3140 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3145 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd279;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3151 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3156 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd280;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd280)) begin
            $error("Failed on action=3161 checking port data_out_data. Expected %x, got %x" , 16'd280, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3162 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3163 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3168 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd281;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3174 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3179 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd282;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd282)) begin
            $error("Failed on action=3184 checking port data_out_data. Expected %x, got %x" , 16'd282, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3185 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3186 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3191 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd283;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3197 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3202 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd284;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd284)) begin
            $error("Failed on action=3207 checking port data_out_data. Expected %x, got %x" , 16'd284, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3208 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3209 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3214 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd285;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3220 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3225 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd286;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd286)) begin
            $error("Failed on action=3230 checking port data_out_data. Expected %x, got %x" , 16'd286, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3231 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3232 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3237 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd287;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3243 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3248 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd288;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3254 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd289;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3265 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd290;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3276 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd291;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3286 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3287 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd292;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3297 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3298 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3303 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd293;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3308 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3309 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3314 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd294;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3319 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3320 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3325 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd295;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3330 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3331 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3336 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd296;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3341 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3342 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3347 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd297;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3352 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3353 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3358 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd298;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3363 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3364 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3369 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd299;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3374 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3375 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3380 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd300;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3385 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3386 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3391 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd301;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3397 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3402 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd302;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3408 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd303;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3419 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd304;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3430 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd305;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3440 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3441 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3446 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd306;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3451 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3452 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3457 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd307;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3462 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3463 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3468 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd308;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3473 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3474 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3479 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd309;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3484 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3485 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3490 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd310;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3495 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3496 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3501 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd311;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3506 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3507 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3512 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd312;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3517 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3518 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3523 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd313;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3528 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3529 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3534 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd314;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3540 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3545 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd315;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3551 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3556 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd316;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3562 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd317;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3573 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd318;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3583 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3584 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3589 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd319;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3594 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3595 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3600 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd320;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd320)) begin
            $error("Failed on action=3605 checking port data_out_data. Expected %x, got %x" , 16'd320, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3606 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3607 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3612 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd321;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3617 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3618 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3623 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd322;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd322)) begin
            $error("Failed on action=3628 checking port data_out_data. Expected %x, got %x" , 16'd322, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3629 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3630 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3635 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd323;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3640 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3641 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3646 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd324;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd324)) begin
            $error("Failed on action=3651 checking port data_out_data. Expected %x, got %x" , 16'd324, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3652 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3653 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3658 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd325;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3663 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3664 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3669 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd326;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd326)) begin
            $error("Failed on action=3674 checking port data_out_data. Expected %x, got %x" , 16'd326, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3675 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3676 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd327;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3686 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3687 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd328;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd328)) begin
            $error("Failed on action=3697 checking port data_out_data. Expected %x, got %x" , 16'd328, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3698 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3699 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd329;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3710 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd330;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd330)) begin
            $error("Failed on action=3720 checking port data_out_data. Expected %x, got %x" , 16'd330, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3721 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3722 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3727 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd331;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3733 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3738 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd332;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd332)) begin
            $error("Failed on action=3743 checking port data_out_data. Expected %x, got %x" , 16'd332, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3744 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3745 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3750 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd333;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3756 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3761 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd334;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd334)) begin
            $error("Failed on action=3766 checking port data_out_data. Expected %x, got %x" , 16'd334, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3767 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3768 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3773 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd335;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3779 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3784 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd336;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd336)) begin
            $error("Failed on action=3789 checking port data_out_data. Expected %x, got %x" , 16'd336, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3790 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3791 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3796 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd337;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3802 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3807 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd338;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd338)) begin
            $error("Failed on action=3812 checking port data_out_data. Expected %x, got %x" , 16'd338, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3813 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3814 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd339;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3825 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd340;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd340)) begin
            $error("Failed on action=3835 checking port data_out_data. Expected %x, got %x" , 16'd340, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3836 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3837 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3842 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd341;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3848 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd342;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd342)) begin
            $error("Failed on action=3858 checking port data_out_data. Expected %x, got %x" , 16'd342, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3859 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3860 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3865 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd343;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3871 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3876 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd344;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd344)) begin
            $error("Failed on action=3881 checking port data_out_data. Expected %x, got %x" , 16'd344, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3882 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3883 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3888 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd345;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3894 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3899 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd346;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd346)) begin
            $error("Failed on action=3904 checking port data_out_data. Expected %x, got %x" , 16'd346, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3905 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3906 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3911 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd347;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3917 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3922 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd348;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd348)) begin
            $error("Failed on action=3927 checking port data_out_data. Expected %x, got %x" , 16'd348, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3928 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3929 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3934 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd349;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3940 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3945 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd350;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd350)) begin
            $error("Failed on action=3950 checking port data_out_data. Expected %x, got %x" , 16'd350, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=3951 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3952 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3957 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd351;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3963 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3968 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd352;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3974 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd353;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3985 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd354;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=3995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=3996 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd355;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4006 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4007 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd356;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4017 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4018 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4023 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd357;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4028 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4029 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4034 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd358;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4039 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4040 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4045 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd359;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4050 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4051 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4056 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd360;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4061 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4062 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4067 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd361;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4072 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4073 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4078 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd362;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4083 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4084 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4089 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd363;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4094 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4095 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4100 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd364;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4105 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4106 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4111 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd365;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4117 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4122 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd366;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4128 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd367;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4139 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4144 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd368;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4149 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4150 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd369;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4160 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4161 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4166 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd370;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4171 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4172 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4177 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd371;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4182 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4183 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4188 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd372;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4193 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4194 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4199 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd373;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4204 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4205 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4210 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd374;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4215 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4216 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4221 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd375;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4226 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4227 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4232 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd376;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4237 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4238 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4243 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd377;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4248 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4249 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4254 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd378;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4260 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4265 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd379;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4271 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd380;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4282 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd381;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4293 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd382;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4303 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4304 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4309 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd383;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4314 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4315 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4320 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd384;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd384)) begin
            $error("Failed on action=4325 checking port data_out_data. Expected %x, got %x" , 16'd384, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4326 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4327 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4332 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd385;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4337 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4338 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4343 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd386;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd386)) begin
            $error("Failed on action=4348 checking port data_out_data. Expected %x, got %x" , 16'd386, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4349 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4350 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4355 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd387;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4360 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4361 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4366 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd388;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd388)) begin
            $error("Failed on action=4371 checking port data_out_data. Expected %x, got %x" , 16'd388, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4372 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4373 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4378 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd389;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4383 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4384 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4389 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd390;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd390)) begin
            $error("Failed on action=4394 checking port data_out_data. Expected %x, got %x" , 16'd390, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4395 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4396 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd391;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4406 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4407 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd392;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd392)) begin
            $error("Failed on action=4417 checking port data_out_data. Expected %x, got %x" , 16'd392, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4418 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4419 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd393;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4430 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd394;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd394)) begin
            $error("Failed on action=4440 checking port data_out_data. Expected %x, got %x" , 16'd394, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4441 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4442 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4447 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd395;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4453 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4458 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd396;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd396)) begin
            $error("Failed on action=4463 checking port data_out_data. Expected %x, got %x" , 16'd396, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4464 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4465 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4470 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd397;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4476 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4481 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd398;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd398)) begin
            $error("Failed on action=4486 checking port data_out_data. Expected %x, got %x" , 16'd398, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4487 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4488 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4493 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd399;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4499 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4504 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd400;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd400)) begin
            $error("Failed on action=4509 checking port data_out_data. Expected %x, got %x" , 16'd400, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4510 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4511 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd401;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4522 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd402;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd402)) begin
            $error("Failed on action=4532 checking port data_out_data. Expected %x, got %x" , 16'd402, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4533 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4534 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd403;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4545 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd404;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd404)) begin
            $error("Failed on action=4555 checking port data_out_data. Expected %x, got %x" , 16'd404, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4556 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4557 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4562 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd405;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4568 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4573 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd406;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd406)) begin
            $error("Failed on action=4578 checking port data_out_data. Expected %x, got %x" , 16'd406, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4579 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4580 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4585 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd407;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4591 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4596 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd408;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd408)) begin
            $error("Failed on action=4601 checking port data_out_data. Expected %x, got %x" , 16'd408, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4602 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4603 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4608 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd409;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4614 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4619 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd410;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd410)) begin
            $error("Failed on action=4624 checking port data_out_data. Expected %x, got %x" , 16'd410, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4625 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4626 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4631 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd411;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4637 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4642 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd412;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd412)) begin
            $error("Failed on action=4647 checking port data_out_data. Expected %x, got %x" , 16'd412, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4648 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4649 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4654 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd413;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4660 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd414;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd414)) begin
            $error("Failed on action=4670 checking port data_out_data. Expected %x, got %x" , 16'd414, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=4671 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4672 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4677 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd415;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4683 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4688 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd416;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4694 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4699 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd417;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4705 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd418;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4716 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4721 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd419;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4726 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4727 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd420;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4737 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4738 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4743 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd421;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4748 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4749 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4754 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd422;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4759 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4760 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4765 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd423;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4770 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4771 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4776 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd424;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4781 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4782 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4787 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd425;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4792 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4793 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4798 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd426;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4803 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4804 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4809 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd427;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4814 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4815 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4820 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd428;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4825 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4826 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4831 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd429;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4837 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4842 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd430;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4848 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd431;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4859 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4864 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd432;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4869 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4870 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd433;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4880 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4881 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4886 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd434;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4891 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4892 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4897 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd435;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4902 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4903 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4908 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd436;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4913 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4914 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4919 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd437;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4924 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4925 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4930 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd438;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4935 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4936 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4941 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd439;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4946 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4947 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4952 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd440;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4957 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4958 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4963 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd441;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4968 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4969 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4974 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd442;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4980 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4985 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd443;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=4991 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=4996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd444;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5002 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd445;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5013 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd446;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5023 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5024 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5029 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd447;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5034 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5035 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5040 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd448;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd448)) begin
            $error("Failed on action=5045 checking port data_out_data. Expected %x, got %x" , 16'd448, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5046 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5047 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5052 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd449;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5057 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5058 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5063 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd450;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd450)) begin
            $error("Failed on action=5068 checking port data_out_data. Expected %x, got %x" , 16'd450, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5069 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5070 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5075 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd451;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5080 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5081 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5086 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd452;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd452)) begin
            $error("Failed on action=5091 checking port data_out_data. Expected %x, got %x" , 16'd452, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5092 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5093 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5098 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd453;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5103 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5104 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5109 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd454;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd454)) begin
            $error("Failed on action=5114 checking port data_out_data. Expected %x, got %x" , 16'd454, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5115 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5116 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd455;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5126 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5127 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd456;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd456)) begin
            $error("Failed on action=5137 checking port data_out_data. Expected %x, got %x" , 16'd456, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5138 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5139 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5144 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd457;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5149 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5150 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd458;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd458)) begin
            $error("Failed on action=5160 checking port data_out_data. Expected %x, got %x" , 16'd458, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5161 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5162 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5167 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd459;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5172 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5173 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5178 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd460;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd460)) begin
            $error("Failed on action=5183 checking port data_out_data. Expected %x, got %x" , 16'd460, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5184 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5185 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5190 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd461;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5195 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5196 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5201 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd462;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd462)) begin
            $error("Failed on action=5206 checking port data_out_data. Expected %x, got %x" , 16'd462, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5207 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5208 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5213 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd463;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5218 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5219 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5224 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd464;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd464)) begin
            $error("Failed on action=5229 checking port data_out_data. Expected %x, got %x" , 16'd464, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5230 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5231 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5236 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd465;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5241 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5242 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd466;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd466)) begin
            $error("Failed on action=5252 checking port data_out_data. Expected %x, got %x" , 16'd466, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5253 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5254 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd467;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5265 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd468;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd468)) begin
            $error("Failed on action=5275 checking port data_out_data. Expected %x, got %x" , 16'd468, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5276 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5277 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5282 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd469;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5288 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5293 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd470;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd470)) begin
            $error("Failed on action=5298 checking port data_out_data. Expected %x, got %x" , 16'd470, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5299 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5300 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5305 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd471;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5310 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5311 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5316 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd472;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd472)) begin
            $error("Failed on action=5321 checking port data_out_data. Expected %x, got %x" , 16'd472, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5322 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5323 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5328 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd473;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5333 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5334 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5339 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd474;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd474)) begin
            $error("Failed on action=5344 checking port data_out_data. Expected %x, got %x" , 16'd474, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5345 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5346 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5351 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd475;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5356 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5357 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5362 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd476;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd476)) begin
            $error("Failed on action=5367 checking port data_out_data. Expected %x, got %x" , 16'd476, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5368 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5369 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5374 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd477;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5380 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5385 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd478;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd478)) begin
            $error("Failed on action=5390 checking port data_out_data. Expected %x, got %x" , 16'd478, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5391 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5392 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5397 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd479;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5402 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5403 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5408 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd480;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5414 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5419 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd481;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5425 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5430 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd482;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5436 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5441 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd483;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5446 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5447 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd484;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5457 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5458 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5463 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd485;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5468 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5469 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5474 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd486;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5479 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5480 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5485 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd487;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5490 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5491 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5496 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd488;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5501 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5502 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5507 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd489;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5512 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5513 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5518 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd490;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5523 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5524 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5529 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd491;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5534 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5535 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5540 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd492;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5545 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5546 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5551 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd493;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5556 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5557 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5562 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd494;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5568 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5573 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd495;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5579 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5584 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd496;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5589 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5590 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5595 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd497;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5600 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5601 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5606 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd498;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5611 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5612 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5617 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd499;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5622 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5623 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5628 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd500;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5633 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5634 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5639 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd501;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5644 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5645 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5650 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd502;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5655 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5656 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5661 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd503;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5666 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5667 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5672 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd504;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5677 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5678 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5683 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd505;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5688 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5689 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5694 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd506;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5699 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5700 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5705 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd507;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5711 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5716 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd508;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5721 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5722 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5727 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd509;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5733 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5738 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd510;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5743 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5744 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5749 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd511;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5754 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5755 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5760 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd512;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd512)) begin
            $error("Failed on action=5765 checking port data_out_data. Expected %x, got %x" , 16'd512, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5766 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5767 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5772 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd513;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5777 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5778 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5783 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd514;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd514)) begin
            $error("Failed on action=5788 checking port data_out_data. Expected %x, got %x" , 16'd514, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5789 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5790 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5795 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd515;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5800 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5801 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5806 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd516;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd516)) begin
            $error("Failed on action=5811 checking port data_out_data. Expected %x, got %x" , 16'd516, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5812 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5813 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5818 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd517;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5823 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5824 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5829 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd518;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd518)) begin
            $error("Failed on action=5834 checking port data_out_data. Expected %x, got %x" , 16'd518, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5835 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5836 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd519;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5846 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5847 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd520;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd520)) begin
            $error("Failed on action=5857 checking port data_out_data. Expected %x, got %x" , 16'd520, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5858 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5859 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5864 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd521;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5869 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5870 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd522;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd522)) begin
            $error("Failed on action=5880 checking port data_out_data. Expected %x, got %x" , 16'd522, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5881 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5882 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5887 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd523;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5892 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5893 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5898 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd524;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd524)) begin
            $error("Failed on action=5903 checking port data_out_data. Expected %x, got %x" , 16'd524, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5904 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5905 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5910 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd525;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5915 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5916 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5921 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd526;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd526)) begin
            $error("Failed on action=5926 checking port data_out_data. Expected %x, got %x" , 16'd526, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5927 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5928 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5933 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd527;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5938 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5939 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5944 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd528;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd528)) begin
            $error("Failed on action=5949 checking port data_out_data. Expected %x, got %x" , 16'd528, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5950 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5951 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5956 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd529;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5961 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5962 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd530;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd530)) begin
            $error("Failed on action=5972 checking port data_out_data. Expected %x, got %x" , 16'd530, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5973 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5974 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd531;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5985 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=5990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd532;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd532)) begin
            $error("Failed on action=5995 checking port data_out_data. Expected %x, got %x" , 16'd532, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=5996 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=5997 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6002 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd533;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6008 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6013 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd534;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd534)) begin
            $error("Failed on action=6018 checking port data_out_data. Expected %x, got %x" , 16'd534, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6019 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6020 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6025 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd535;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6030 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6031 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6036 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd536;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd536)) begin
            $error("Failed on action=6041 checking port data_out_data. Expected %x, got %x" , 16'd536, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6042 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6043 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6048 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd537;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6053 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6054 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6059 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd538;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd538)) begin
            $error("Failed on action=6064 checking port data_out_data. Expected %x, got %x" , 16'd538, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6065 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6066 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6071 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd539;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6076 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6077 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6082 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd540;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd540)) begin
            $error("Failed on action=6087 checking port data_out_data. Expected %x, got %x" , 16'd540, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6088 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6089 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6094 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd541;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6100 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6105 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd542;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd542)) begin
            $error("Failed on action=6110 checking port data_out_data. Expected %x, got %x" , 16'd542, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6111 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6112 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6117 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd543;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6122 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6123 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6128 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd544;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6134 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6139 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd545;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6144 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6145 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd546;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6156 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6161 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd547;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6166 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6167 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6172 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd548;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6177 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6178 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6183 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd549;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6188 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6189 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6194 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd550;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6199 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6200 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6205 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd551;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6210 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6211 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6216 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd552;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6221 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6222 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6227 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd553;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6232 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6233 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6238 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd554;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6243 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6244 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6249 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd555;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6254 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6255 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6260 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd556;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6265 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6266 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6271 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd557;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6277 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6282 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd558;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6288 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6293 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd559;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6299 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6304 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd560;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6309 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6310 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6315 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd561;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6320 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6321 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6326 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd562;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6331 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6332 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6337 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd563;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6342 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6343 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6348 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd564;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6353 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6354 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6359 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd565;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6364 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6365 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6370 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd566;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6375 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6376 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6381 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd567;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6386 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6387 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6392 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd568;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6397 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6398 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6403 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd569;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6408 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6409 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6414 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd570;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6419 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6420 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6425 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd571;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6430 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6431 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6436 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd572;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6441 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6442 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6447 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd573;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6453 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6458 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd574;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6463 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6464 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6469 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd575;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6474 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6475 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6480 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd576;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd576)) begin
            $error("Failed on action=6485 checking port data_out_data. Expected %x, got %x" , 16'd576, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6486 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6487 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6492 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd577;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6497 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6498 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6503 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd578;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd578)) begin
            $error("Failed on action=6508 checking port data_out_data. Expected %x, got %x" , 16'd578, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6509 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6510 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6515 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd579;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6520 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6521 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6526 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd580;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd580)) begin
            $error("Failed on action=6531 checking port data_out_data. Expected %x, got %x" , 16'd580, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6532 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6533 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6538 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd581;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6543 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6544 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6549 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd582;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd582)) begin
            $error("Failed on action=6554 checking port data_out_data. Expected %x, got %x" , 16'd582, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6555 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6556 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd583;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6566 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6567 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd584;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd584)) begin
            $error("Failed on action=6577 checking port data_out_data. Expected %x, got %x" , 16'd584, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6578 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6579 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6584 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd585;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6589 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6590 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6595 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd586;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd586)) begin
            $error("Failed on action=6600 checking port data_out_data. Expected %x, got %x" , 16'd586, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6601 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6602 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6607 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd587;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6612 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6613 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6618 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd588;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd588)) begin
            $error("Failed on action=6623 checking port data_out_data. Expected %x, got %x" , 16'd588, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6624 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6625 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6630 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd589;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6635 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6636 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6641 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd590;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd590)) begin
            $error("Failed on action=6646 checking port data_out_data. Expected %x, got %x" , 16'd590, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6647 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6648 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6653 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd591;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6658 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6659 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6664 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd592;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd592)) begin
            $error("Failed on action=6669 checking port data_out_data. Expected %x, got %x" , 16'd592, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6670 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6671 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd593;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6682 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd594;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd594)) begin
            $error("Failed on action=6692 checking port data_out_data. Expected %x, got %x" , 16'd594, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6693 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6694 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6699 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd595;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6705 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd596;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd596)) begin
            $error("Failed on action=6715 checking port data_out_data. Expected %x, got %x" , 16'd596, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6716 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6717 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6722 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd597;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6727 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6728 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6733 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd598;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd598)) begin
            $error("Failed on action=6738 checking port data_out_data. Expected %x, got %x" , 16'd598, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6739 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6740 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6745 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd599;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6750 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6751 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6756 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd600;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd600)) begin
            $error("Failed on action=6761 checking port data_out_data. Expected %x, got %x" , 16'd600, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6762 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6763 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6768 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd601;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6773 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6774 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6779 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd602;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd602)) begin
            $error("Failed on action=6784 checking port data_out_data. Expected %x, got %x" , 16'd602, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6785 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6786 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6791 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd603;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6796 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6797 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6802 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd604;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd604)) begin
            $error("Failed on action=6807 checking port data_out_data. Expected %x, got %x" , 16'd604, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6808 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6809 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6814 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd605;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6820 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6825 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd606;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd606)) begin
            $error("Failed on action=6830 checking port data_out_data. Expected %x, got %x" , 16'd606, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=6831 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6832 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6837 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd607;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6842 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6843 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6848 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd608;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6854 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6859 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd609;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6864 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6865 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd610;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6876 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6881 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd611;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6886 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6887 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6892 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd612;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6897 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6898 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6903 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd613;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6908 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6909 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6914 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd614;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6919 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6920 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6925 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd615;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6930 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6931 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6936 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd616;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6941 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6942 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6947 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd617;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6952 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6953 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6958 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd618;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6963 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6964 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6969 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd619;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6974 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6975 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6980 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd620;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6985 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6986 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6991 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd621;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=6996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=6997 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7002 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd622;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7008 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7013 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd623;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7019 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7024 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd624;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7029 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7030 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7035 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd625;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7040 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7041 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7046 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd626;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7051 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7052 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7057 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd627;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7062 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7063 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7068 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd628;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7073 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7074 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7079 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd629;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7084 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7085 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7090 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd630;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7095 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7096 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7101 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd631;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7106 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7107 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7112 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd632;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7117 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7118 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7123 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd633;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7128 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7129 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7134 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd634;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7139 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7140 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7145 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd635;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7151 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7156 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd636;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7161 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7162 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7167 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd637;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7172 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7173 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7178 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd638;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7183 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7184 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7189 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd639;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7194 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7195 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7200 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd640;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd640)) begin
            $error("Failed on action=7205 checking port data_out_data. Expected %x, got %x" , 16'd640, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7206 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7207 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7212 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd641;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7217 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7218 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7223 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd642;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd642)) begin
            $error("Failed on action=7228 checking port data_out_data. Expected %x, got %x" , 16'd642, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7229 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7230 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7235 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd643;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7240 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7241 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7246 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd644;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd644)) begin
            $error("Failed on action=7251 checking port data_out_data. Expected %x, got %x" , 16'd644, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7252 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7253 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7258 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd645;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7263 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7264 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7269 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd646;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd646)) begin
            $error("Failed on action=7274 checking port data_out_data. Expected %x, got %x" , 16'd646, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7275 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7276 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd647;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7286 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7287 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd648;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd648)) begin
            $error("Failed on action=7297 checking port data_out_data. Expected %x, got %x" , 16'd648, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7298 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7299 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7304 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd649;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7309 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7310 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7315 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd650;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd650)) begin
            $error("Failed on action=7320 checking port data_out_data. Expected %x, got %x" , 16'd650, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7321 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7322 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7327 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd651;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7332 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7333 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7338 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd652;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd652)) begin
            $error("Failed on action=7343 checking port data_out_data. Expected %x, got %x" , 16'd652, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7344 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7345 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7350 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd653;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7355 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7356 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7361 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd654;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd654)) begin
            $error("Failed on action=7366 checking port data_out_data. Expected %x, got %x" , 16'd654, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7367 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7368 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7373 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd655;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7378 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7379 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd656;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd656)) begin
            $error("Failed on action=7389 checking port data_out_data. Expected %x, got %x" , 16'd656, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7390 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7391 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd657;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7402 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd658;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd658)) begin
            $error("Failed on action=7412 checking port data_out_data. Expected %x, got %x" , 16'd658, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7413 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7414 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7419 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd659;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7425 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7430 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd660;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd660)) begin
            $error("Failed on action=7435 checking port data_out_data. Expected %x, got %x" , 16'd660, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7436 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7437 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7442 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd661;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7447 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7448 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7453 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd662;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd662)) begin
            $error("Failed on action=7458 checking port data_out_data. Expected %x, got %x" , 16'd662, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7459 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7460 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7465 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd663;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7470 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7471 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7476 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd664;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd664)) begin
            $error("Failed on action=7481 checking port data_out_data. Expected %x, got %x" , 16'd664, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7482 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7483 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7488 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd665;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7493 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7494 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7499 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd666;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd666)) begin
            $error("Failed on action=7504 checking port data_out_data. Expected %x, got %x" , 16'd666, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7505 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7506 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7511 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd667;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7517 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7522 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd668;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd668)) begin
            $error("Failed on action=7527 checking port data_out_data. Expected %x, got %x" , 16'd668, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7528 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7529 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7534 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd669;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7540 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7545 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd670;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd670)) begin
            $error("Failed on action=7550 checking port data_out_data. Expected %x, got %x" , 16'd670, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7551 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7552 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7557 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd671;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7562 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7563 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7568 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd672;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7573 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7574 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7579 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd673;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7584 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7585 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd674;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7595 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7596 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7601 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd675;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7606 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7607 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7612 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd676;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7617 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7618 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7623 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd677;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7628 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7629 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7634 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd678;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7639 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7640 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7645 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd679;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7650 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7651 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7656 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd680;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7661 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7662 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7667 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd681;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7672 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7673 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7678 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd682;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7683 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7684 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7689 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd683;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7694 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7695 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7700 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd684;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7705 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7706 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7711 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd685;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7716 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7717 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7722 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd686;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7727 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7728 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7733 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd687;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7738 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7739 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7744 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd688;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7749 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7750 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd689;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7760 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7761 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7766 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd690;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7771 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7772 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7777 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd691;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7782 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7783 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7788 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd692;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7793 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7794 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7799 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd693;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7804 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7805 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7810 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd694;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7815 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7816 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7821 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd695;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7826 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7827 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7832 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd696;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7837 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7838 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7843 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd697;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7848 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7849 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7854 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd698;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7859 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7860 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7865 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd699;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7871 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7876 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd700;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7881 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7882 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7887 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd701;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7892 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7893 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7898 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd702;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7903 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7904 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7909 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd703;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7914 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7915 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7920 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd704;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd704)) begin
            $error("Failed on action=7925 checking port data_out_data. Expected %x, got %x" , 16'd704, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7926 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7927 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7932 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd705;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7937 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7938 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7943 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd706;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd706)) begin
            $error("Failed on action=7948 checking port data_out_data. Expected %x, got %x" , 16'd706, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7949 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7950 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7955 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd707;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7960 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7961 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7966 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd708;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd708)) begin
            $error("Failed on action=7971 checking port data_out_data. Expected %x, got %x" , 16'd708, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7972 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7973 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7978 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd709;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7983 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7984 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=7989 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd710;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd710)) begin
            $error("Failed on action=7994 checking port data_out_data. Expected %x, got %x" , 16'd710, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=7995 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=7996 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd711;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8006 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8007 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd712;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd712)) begin
            $error("Failed on action=8017 checking port data_out_data. Expected %x, got %x" , 16'd712, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8018 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8019 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8024 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd713;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8029 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8030 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8035 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd714;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd714)) begin
            $error("Failed on action=8040 checking port data_out_data. Expected %x, got %x" , 16'd714, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8041 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8042 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8047 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd715;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8052 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8053 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8058 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd716;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd716)) begin
            $error("Failed on action=8063 checking port data_out_data. Expected %x, got %x" , 16'd716, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8064 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8065 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8070 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd717;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8075 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8076 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8081 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd718;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd718)) begin
            $error("Failed on action=8086 checking port data_out_data. Expected %x, got %x" , 16'd718, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8087 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8088 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8093 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd719;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8098 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8099 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd720;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd720)) begin
            $error("Failed on action=8109 checking port data_out_data. Expected %x, got %x" , 16'd720, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8110 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8111 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd721;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8122 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd722;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd722)) begin
            $error("Failed on action=8132 checking port data_out_data. Expected %x, got %x" , 16'd722, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8133 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8134 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8139 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd723;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8144 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8145 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd724;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd724)) begin
            $error("Failed on action=8155 checking port data_out_data. Expected %x, got %x" , 16'd724, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8156 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8157 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8162 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd725;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8167 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8168 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd726;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd726)) begin
            $error("Failed on action=8178 checking port data_out_data. Expected %x, got %x" , 16'd726, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8179 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8180 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8185 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd727;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8190 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8191 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd728;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd728)) begin
            $error("Failed on action=8201 checking port data_out_data. Expected %x, got %x" , 16'd728, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8202 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8203 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8208 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd729;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8213 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8214 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd730;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd730)) begin
            $error("Failed on action=8224 checking port data_out_data. Expected %x, got %x" , 16'd730, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8225 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8226 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8231 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd731;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8236 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8237 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd732;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd732)) begin
            $error("Failed on action=8247 checking port data_out_data. Expected %x, got %x" , 16'd732, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8248 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8249 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8254 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd733;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8260 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8265 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd734;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd734)) begin
            $error("Failed on action=8270 checking port data_out_data. Expected %x, got %x" , 16'd734, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8271 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8272 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8277 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd735;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8282 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8283 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8288 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd736;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8293 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8294 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8299 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd737;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8304 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8305 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8310 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd738;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8315 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8316 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8321 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd739;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8326 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8327 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8332 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd740;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8337 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8338 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8343 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd741;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8348 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8349 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8354 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd742;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8359 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8360 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8365 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd743;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8370 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8371 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8376 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd744;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8381 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8382 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8387 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd745;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8392 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8393 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8398 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd746;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8403 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8404 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8409 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd747;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8414 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8415 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8420 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd748;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8425 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8426 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8431 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd749;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8436 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8437 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8442 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd750;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8447 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8448 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8453 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd751;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8458 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8459 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8464 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd752;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8469 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8470 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd753;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8480 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8481 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8486 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd754;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8491 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8492 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8497 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd755;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8502 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8503 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8508 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd756;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8513 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8514 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8519 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd757;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8524 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8525 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8530 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd758;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8535 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8536 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8541 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd759;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8546 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8547 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8552 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd760;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8557 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8558 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8563 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd761;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8568 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8569 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8574 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd762;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8579 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8580 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8585 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd763;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8591 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8596 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd764;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8601 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8602 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8607 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd765;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8612 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8613 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8618 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd766;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8623 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8624 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8629 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd767;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8634 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8635 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8640 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd768;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd768)) begin
            $error("Failed on action=8645 checking port data_out_data. Expected %x, got %x" , 16'd768, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8646 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8647 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8652 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd769;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8657 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8658 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8663 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd770;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd770)) begin
            $error("Failed on action=8668 checking port data_out_data. Expected %x, got %x" , 16'd770, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8669 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8670 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8675 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd771;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8680 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8681 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8686 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd772;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd772)) begin
            $error("Failed on action=8691 checking port data_out_data. Expected %x, got %x" , 16'd772, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8692 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8693 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd773;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8703 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8704 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd774;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd774)) begin
            $error("Failed on action=8714 checking port data_out_data. Expected %x, got %x" , 16'd774, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8715 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8716 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8721 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd775;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8726 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8727 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd776;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd776)) begin
            $error("Failed on action=8737 checking port data_out_data. Expected %x, got %x" , 16'd776, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8738 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8739 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8744 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd777;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8749 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8750 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd778;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd778)) begin
            $error("Failed on action=8760 checking port data_out_data. Expected %x, got %x" , 16'd778, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8761 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8762 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8767 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd779;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8772 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8773 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd780;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd780)) begin
            $error("Failed on action=8783 checking port data_out_data. Expected %x, got %x" , 16'd780, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8784 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8785 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8790 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd781;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8795 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8796 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd782;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd782)) begin
            $error("Failed on action=8806 checking port data_out_data. Expected %x, got %x" , 16'd782, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8807 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8808 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8813 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd783;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8818 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8819 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd784;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd784)) begin
            $error("Failed on action=8829 checking port data_out_data. Expected %x, got %x" , 16'd784, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8830 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8831 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd785;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8842 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd786;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd786)) begin
            $error("Failed on action=8852 checking port data_out_data. Expected %x, got %x" , 16'd786, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8853 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8854 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8859 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd787;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8864 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8865 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd788;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd788)) begin
            $error("Failed on action=8875 checking port data_out_data. Expected %x, got %x" , 16'd788, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8876 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8877 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8882 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd789;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8887 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8888 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd790;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd790)) begin
            $error("Failed on action=8898 checking port data_out_data. Expected %x, got %x" , 16'd790, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8899 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8900 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8905 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd791;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8910 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8911 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd792;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd792)) begin
            $error("Failed on action=8921 checking port data_out_data. Expected %x, got %x" , 16'd792, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8922 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8923 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8928 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd793;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8933 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8934 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd794;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd794)) begin
            $error("Failed on action=8944 checking port data_out_data. Expected %x, got %x" , 16'd794, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8945 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8946 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8951 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd795;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8956 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8957 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd796;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd796)) begin
            $error("Failed on action=8967 checking port data_out_data. Expected %x, got %x" , 16'd796, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8968 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8969 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8974 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd797;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8980 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8985 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd798;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd798)) begin
            $error("Failed on action=8990 checking port data_out_data. Expected %x, got %x" , 16'd798, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=8991 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=8992 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=8997 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd799;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9002 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9003 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9008 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd800;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9013 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9014 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9019 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd801;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9024 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9025 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9030 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd802;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9035 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9036 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9041 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd803;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9046 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9047 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9052 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd804;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9057 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9058 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9063 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd805;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9068 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9069 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9074 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd806;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9079 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9080 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9085 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd807;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9090 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9091 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9096 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd808;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9101 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9102 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9107 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd809;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9112 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9113 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9118 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd810;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9123 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9124 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9129 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd811;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9134 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9135 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9140 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd812;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9145 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9146 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9151 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd813;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9156 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9157 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9162 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd814;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9167 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9168 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd815;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9178 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9179 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9184 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd816;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9189 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9190 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9195 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd817;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9200 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9201 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9206 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd818;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9211 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9212 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9217 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd819;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9222 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9223 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9228 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd820;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9233 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9234 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9239 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd821;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9244 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9245 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9250 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd822;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9255 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9256 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9261 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd823;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9266 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9267 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9272 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd824;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9277 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9278 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9283 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd825;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9288 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9289 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9294 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd826;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9299 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9300 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9305 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd827;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9310 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9311 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9316 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd828;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9321 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9322 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9327 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd829;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9332 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9333 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9338 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd830;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9343 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9344 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9349 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd831;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9354 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9355 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9360 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd832;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd832)) begin
            $error("Failed on action=9365 checking port data_out_data. Expected %x, got %x" , 16'd832, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9366 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9367 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9372 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd833;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9377 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9378 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9383 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd834;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd834)) begin
            $error("Failed on action=9388 checking port data_out_data. Expected %x, got %x" , 16'd834, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9389 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9390 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9395 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd835;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9400 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9401 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9406 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd836;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd836)) begin
            $error("Failed on action=9411 checking port data_out_data. Expected %x, got %x" , 16'd836, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9412 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9413 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd837;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9423 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9424 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd838;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd838)) begin
            $error("Failed on action=9434 checking port data_out_data. Expected %x, got %x" , 16'd838, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9435 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9436 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9441 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd839;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9446 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9447 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd840;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd840)) begin
            $error("Failed on action=9457 checking port data_out_data. Expected %x, got %x" , 16'd840, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9458 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9459 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9464 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd841;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9469 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9470 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd842;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd842)) begin
            $error("Failed on action=9480 checking port data_out_data. Expected %x, got %x" , 16'd842, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9481 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9482 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9487 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd843;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9492 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9493 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd844;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd844)) begin
            $error("Failed on action=9503 checking port data_out_data. Expected %x, got %x" , 16'd844, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9504 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9505 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9510 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd845;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9515 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9516 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd846;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd846)) begin
            $error("Failed on action=9526 checking port data_out_data. Expected %x, got %x" , 16'd846, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9527 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9528 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd847;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9538 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9539 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd848;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd848)) begin
            $error("Failed on action=9549 checking port data_out_data. Expected %x, got %x" , 16'd848, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9550 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9551 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9556 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd849;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9562 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd850;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd850)) begin
            $error("Failed on action=9572 checking port data_out_data. Expected %x, got %x" , 16'd850, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9573 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9574 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9579 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd851;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9584 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9585 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd852;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd852)) begin
            $error("Failed on action=9595 checking port data_out_data. Expected %x, got %x" , 16'd852, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9596 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9597 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9602 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd853;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9607 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9608 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd854;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd854)) begin
            $error("Failed on action=9618 checking port data_out_data. Expected %x, got %x" , 16'd854, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9619 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9620 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9625 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd855;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9630 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9631 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd856;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd856)) begin
            $error("Failed on action=9641 checking port data_out_data. Expected %x, got %x" , 16'd856, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9642 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9643 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9648 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd857;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9653 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9654 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd858;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd858)) begin
            $error("Failed on action=9664 checking port data_out_data. Expected %x, got %x" , 16'd858, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9665 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9666 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9671 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd859;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9677 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd860;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd860)) begin
            $error("Failed on action=9687 checking port data_out_data. Expected %x, got %x" , 16'd860, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9688 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9689 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9694 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd861;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9699 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9700 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9705 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd862;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd862)) begin
            $error("Failed on action=9710 checking port data_out_data. Expected %x, got %x" , 16'd862, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=9711 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9712 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9717 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd863;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9722 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9723 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9728 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd864;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9733 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9734 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9739 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd865;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9744 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9745 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9750 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd866;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9756 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9761 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd867;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9766 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9767 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9772 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd868;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9777 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9778 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9783 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd869;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9788 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9789 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9794 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd870;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9799 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9800 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9805 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd871;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9810 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9811 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9816 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd872;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9821 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9822 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9827 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd873;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9832 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9833 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9838 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd874;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9843 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9844 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9849 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd875;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9854 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9855 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9860 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd876;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9865 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9866 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9871 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd877;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9876 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9877 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9882 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd878;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9887 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9888 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd879;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9898 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9899 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9904 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd880;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9909 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9910 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9915 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd881;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9920 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9921 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9926 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd882;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9931 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9932 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9937 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd883;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9942 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9943 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9948 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd884;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9953 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9954 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9959 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd885;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9964 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9965 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9970 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd886;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9975 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9976 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9981 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd887;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9986 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9987 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9992 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd888;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=9997 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=9998 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10003 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd889;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10008 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10009 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10014 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd890;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10019 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10020 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10025 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd891;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10030 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10031 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10036 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd892;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10041 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10042 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10047 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd893;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10052 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10053 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10058 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd894;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10063 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10064 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10069 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd895;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10074 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10075 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10080 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd896;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd896)) begin
            $error("Failed on action=10085 checking port data_out_data. Expected %x, got %x" , 16'd896, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10086 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10087 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10092 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd897;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10097 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10098 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10103 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd898;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd898)) begin
            $error("Failed on action=10108 checking port data_out_data. Expected %x, got %x" , 16'd898, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10109 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10110 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd899;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10120 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10121 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10126 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd900;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd900)) begin
            $error("Failed on action=10131 checking port data_out_data. Expected %x, got %x" , 16'd900, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10132 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10133 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd901;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10143 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10144 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10149 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd902;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd902)) begin
            $error("Failed on action=10154 checking port data_out_data. Expected %x, got %x" , 16'd902, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10155 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10156 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10161 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd903;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10166 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10167 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10172 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd904;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd904)) begin
            $error("Failed on action=10177 checking port data_out_data. Expected %x, got %x" , 16'd904, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10178 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10179 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10184 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd905;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10189 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10190 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10195 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd906;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd906)) begin
            $error("Failed on action=10200 checking port data_out_data. Expected %x, got %x" , 16'd906, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10201 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10202 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10207 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd907;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10212 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10213 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10218 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd908;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd908)) begin
            $error("Failed on action=10223 checking port data_out_data. Expected %x, got %x" , 16'd908, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10224 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10225 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10230 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd909;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10235 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10236 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10241 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd910;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd910)) begin
            $error("Failed on action=10246 checking port data_out_data. Expected %x, got %x" , 16'd910, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10247 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10248 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd911;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10258 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10259 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd912;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd912)) begin
            $error("Failed on action=10269 checking port data_out_data. Expected %x, got %x" , 16'd912, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10270 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10271 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd913;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10282 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd914;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd914)) begin
            $error("Failed on action=10292 checking port data_out_data. Expected %x, got %x" , 16'd914, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10293 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10294 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10299 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd915;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10304 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10305 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10310 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd916;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd916)) begin
            $error("Failed on action=10315 checking port data_out_data. Expected %x, got %x" , 16'd916, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10316 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10317 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10322 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd917;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10327 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10328 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10333 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd918;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd918)) begin
            $error("Failed on action=10338 checking port data_out_data. Expected %x, got %x" , 16'd918, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10339 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10340 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10345 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd919;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10350 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10351 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10356 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd920;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd920)) begin
            $error("Failed on action=10361 checking port data_out_data. Expected %x, got %x" , 16'd920, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10362 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10363 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10368 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd921;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10373 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10374 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd922;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd922)) begin
            $error("Failed on action=10384 checking port data_out_data. Expected %x, got %x" , 16'd922, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10385 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10386 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10391 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd923;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10397 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10402 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd924;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd924)) begin
            $error("Failed on action=10407 checking port data_out_data. Expected %x, got %x" , 16'd924, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10408 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10409 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10414 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd925;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10419 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10420 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10425 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd926;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd926)) begin
            $error("Failed on action=10430 checking port data_out_data. Expected %x, got %x" , 16'd926, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10431 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10432 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10437 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd927;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10442 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10443 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10448 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd928;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10453 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10454 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10459 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd929;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10464 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10465 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10470 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd930;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10476 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10481 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd931;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10486 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10487 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10492 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd932;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10497 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10498 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10503 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd933;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10508 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10509 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10514 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd934;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10519 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10520 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10525 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd935;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10530 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10531 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10536 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd936;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10541 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10542 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10547 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd937;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10552 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10553 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10558 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd938;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10563 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10564 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10569 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd939;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10574 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10575 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10580 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd940;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10585 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10586 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10591 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd941;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10596 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10597 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10602 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd942;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10607 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10608 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd943;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10618 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10619 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10624 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd944;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10629 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10630 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10635 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd945;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10640 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10641 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10646 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd946;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10651 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10652 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10657 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd947;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10662 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10663 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10668 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd948;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10673 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10674 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10679 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd949;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10684 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10685 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10690 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd950;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10695 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10696 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10701 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd951;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10706 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10707 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10712 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd952;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10717 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10718 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10723 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd953;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10728 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10729 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10734 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd954;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10739 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10740 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10745 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd955;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10750 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10751 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10756 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd956;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10761 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10762 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10767 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd957;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10772 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10773 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd958;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10783 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10784 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10789 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd959;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10794 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10795 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10800 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd960;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd960)) begin
            $error("Failed on action=10805 checking port data_out_data. Expected %x, got %x" , 16'd960, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10806 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10807 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10812 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd961;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10817 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10818 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10823 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd962;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd962)) begin
            $error("Failed on action=10828 checking port data_out_data. Expected %x, got %x" , 16'd962, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10829 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10830 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd963;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10840 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10841 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10846 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd964;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd964)) begin
            $error("Failed on action=10851 checking port data_out_data. Expected %x, got %x" , 16'd964, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10852 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10853 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd965;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10863 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10864 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10869 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd966;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd966)) begin
            $error("Failed on action=10874 checking port data_out_data. Expected %x, got %x" , 16'd966, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10875 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10876 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10881 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd967;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10886 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10887 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10892 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd968;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd968)) begin
            $error("Failed on action=10897 checking port data_out_data. Expected %x, got %x" , 16'd968, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10898 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10899 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10904 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd969;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10909 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10910 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10915 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd970;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd970)) begin
            $error("Failed on action=10920 checking port data_out_data. Expected %x, got %x" , 16'd970, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10921 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10922 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10927 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd971;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10932 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10933 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10938 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd972;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd972)) begin
            $error("Failed on action=10943 checking port data_out_data. Expected %x, got %x" , 16'd972, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10944 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10945 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10950 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd973;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10955 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10956 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10961 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd974;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd974)) begin
            $error("Failed on action=10966 checking port data_out_data. Expected %x, got %x" , 16'd974, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10967 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10968 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd975;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10978 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10979 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd976;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd976)) begin
            $error("Failed on action=10989 checking port data_out_data. Expected %x, got %x" , 16'd976, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=10990 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=10991 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=10996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd977;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11002 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd978;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd978)) begin
            $error("Failed on action=11012 checking port data_out_data. Expected %x, got %x" , 16'd978, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11013 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11014 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11019 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd979;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11024 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11025 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11030 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd980;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd980)) begin
            $error("Failed on action=11035 checking port data_out_data. Expected %x, got %x" , 16'd980, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11036 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11037 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11042 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd981;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11047 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11048 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11053 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd982;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd982)) begin
            $error("Failed on action=11058 checking port data_out_data. Expected %x, got %x" , 16'd982, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11059 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11060 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11065 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd983;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11070 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11071 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11076 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd984;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd984)) begin
            $error("Failed on action=11081 checking port data_out_data. Expected %x, got %x" , 16'd984, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11082 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11083 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11088 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd985;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11093 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11094 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd986;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd986)) begin
            $error("Failed on action=11104 checking port data_out_data. Expected %x, got %x" , 16'd986, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11105 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11106 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11111 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd987;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11117 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11122 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd988;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd988)) begin
            $error("Failed on action=11127 checking port data_out_data. Expected %x, got %x" , 16'd988, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11128 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11129 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11134 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd989;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11139 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11140 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11145 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd990;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd990)) begin
            $error("Failed on action=11150 checking port data_out_data. Expected %x, got %x" , 16'd990, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11151 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11152 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11157 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd991;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11162 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11163 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11168 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd992;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11174 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11179 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd993;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11184 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11185 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11190 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd994;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11195 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11196 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11201 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd995;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11206 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11207 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11212 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd996;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11217 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11218 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11223 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd997;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11228 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11229 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11234 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd998;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11239 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11240 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11245 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd999;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11250 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11251 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11256 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1000;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11261 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11262 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11267 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1001;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11272 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11273 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11278 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1002;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11283 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11284 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11289 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1003;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11294 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11295 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11300 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1004;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11305 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11306 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11311 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1005;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11316 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11317 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11322 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1006;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11327 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11328 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11333 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1007;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11338 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11339 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11344 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1008;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11349 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11350 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11355 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1009;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11360 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11361 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11366 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1010;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11371 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11372 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11377 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1011;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11382 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11383 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11388 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1012;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11393 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11394 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11399 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1013;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11404 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11405 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11410 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1014;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11415 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11416 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11421 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1015;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11426 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11427 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11432 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1016;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11437 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11438 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11443 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1017;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11448 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11449 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11454 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1018;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11459 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11460 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11465 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1019;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11470 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11471 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11476 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1020;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11481 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11482 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11487 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1021;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11492 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11493 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1022;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11503 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11504 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11509 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1023;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11514 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11515 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11520 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd0;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd0)) begin
            $error("Failed on action=11525 checking port data_out_data. Expected %x, got %x" , 16'd0, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11526 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11527 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11532 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11537 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11538 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11543 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd2;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd2)) begin
            $error("Failed on action=11548 checking port data_out_data. Expected %x, got %x" , 16'd2, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11549 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11550 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd3;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11560 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11561 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11566 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd4;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd4)) begin
            $error("Failed on action=11571 checking port data_out_data. Expected %x, got %x" , 16'd4, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11572 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11573 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd5;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11583 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11584 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11589 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd6;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd6)) begin
            $error("Failed on action=11594 checking port data_out_data. Expected %x, got %x" , 16'd6, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11595 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11596 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11601 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd7;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11606 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11607 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11612 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd8;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd8)) begin
            $error("Failed on action=11617 checking port data_out_data. Expected %x, got %x" , 16'd8, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11618 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11619 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11624 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd9;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11629 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11630 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11635 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd10;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd10)) begin
            $error("Failed on action=11640 checking port data_out_data. Expected %x, got %x" , 16'd10, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11641 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11642 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11647 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd11;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11652 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11653 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11658 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd12;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd12)) begin
            $error("Failed on action=11663 checking port data_out_data. Expected %x, got %x" , 16'd12, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11664 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11665 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd13;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11675 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11676 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd14;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd14)) begin
            $error("Failed on action=11686 checking port data_out_data. Expected %x, got %x" , 16'd14, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11687 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11688 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd15;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11699 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd16;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd16)) begin
            $error("Failed on action=11709 checking port data_out_data. Expected %x, got %x" , 16'd16, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11710 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11711 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11716 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd17;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11721 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11722 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11727 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd18;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd18)) begin
            $error("Failed on action=11732 checking port data_out_data. Expected %x, got %x" , 16'd18, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11733 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11734 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11739 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd19;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11744 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11745 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11750 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd20;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd20)) begin
            $error("Failed on action=11755 checking port data_out_data. Expected %x, got %x" , 16'd20, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11756 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11757 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11762 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd21;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11767 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11768 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11773 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd22;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd22)) begin
            $error("Failed on action=11778 checking port data_out_data. Expected %x, got %x" , 16'd22, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11779 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11780 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11785 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd23;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11790 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11791 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11796 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd24;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd24)) begin
            $error("Failed on action=11801 checking port data_out_data. Expected %x, got %x" , 16'd24, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11802 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11803 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11808 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd25;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11813 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11814 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd26;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd26)) begin
            $error("Failed on action=11824 checking port data_out_data. Expected %x, got %x" , 16'd26, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11825 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11826 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11831 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd27;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11837 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11842 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd28;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd28)) begin
            $error("Failed on action=11847 checking port data_out_data. Expected %x, got %x" , 16'd28, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11848 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11849 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11854 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd29;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11859 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11860 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11865 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd30;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd30)) begin
            $error("Failed on action=11870 checking port data_out_data. Expected %x, got %x" , 16'd30, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=11871 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11872 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11877 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd31;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11882 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11883 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11888 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd32;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11894 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11899 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd33;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11904 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11905 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11910 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd34;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11915 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11916 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11921 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd35;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11926 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11927 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11932 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd36;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11937 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11938 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11943 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd37;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11948 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11949 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11954 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd38;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11959 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11960 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11965 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd39;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11970 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11971 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11976 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd40;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11981 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11982 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11987 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd41;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11992 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=11993 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=11998 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd42;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12003 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12004 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12009 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd43;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12014 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12015 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12020 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd44;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12025 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12026 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12031 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd45;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12036 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12037 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12042 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd46;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12047 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12048 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12053 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd47;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12058 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12059 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12064 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd48;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12069 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12070 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12075 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd49;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12080 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12081 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12086 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd50;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12091 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12092 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12097 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd51;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12102 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12103 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12108 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd52;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12113 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12114 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12119 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd53;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12124 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12125 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12130 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd54;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12135 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12136 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12141 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd55;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12146 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12147 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12152 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd56;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12157 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12158 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12163 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd57;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12168 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12169 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12174 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd58;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12179 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12180 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12185 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd59;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12190 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12191 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd60;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12201 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12202 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12207 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd61;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12212 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12213 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12218 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd62;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12223 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12224 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12229 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd63;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12234 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12235 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12240 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd64;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd64)) begin
            $error("Failed on action=12245 checking port data_out_data. Expected %x, got %x" , 16'd64, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12246 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12247 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12252 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd65;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12257 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12258 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12263 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd66;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd66)) begin
            $error("Failed on action=12268 checking port data_out_data. Expected %x, got %x" , 16'd66, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12269 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12270 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd67;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12280 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12281 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12286 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd68;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd68)) begin
            $error("Failed on action=12291 checking port data_out_data. Expected %x, got %x" , 16'd68, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12292 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12293 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd69;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12303 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12304 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12309 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd70;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd70)) begin
            $error("Failed on action=12314 checking port data_out_data. Expected %x, got %x" , 16'd70, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12315 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12316 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12321 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd71;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12326 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12327 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12332 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd72;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd72)) begin
            $error("Failed on action=12337 checking port data_out_data. Expected %x, got %x" , 16'd72, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12338 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12339 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12344 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd73;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12349 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12350 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12355 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd74;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd74)) begin
            $error("Failed on action=12360 checking port data_out_data. Expected %x, got %x" , 16'd74, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12361 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12362 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12367 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd75;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12372 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12373 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12378 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd76;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd76)) begin
            $error("Failed on action=12383 checking port data_out_data. Expected %x, got %x" , 16'd76, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12384 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12385 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd77;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12395 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12396 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd78;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd78)) begin
            $error("Failed on action=12406 checking port data_out_data. Expected %x, got %x" , 16'd78, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12407 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12408 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd79;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12419 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd80;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd80)) begin
            $error("Failed on action=12429 checking port data_out_data. Expected %x, got %x" , 16'd80, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12430 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12431 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12436 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd81;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12441 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12442 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12447 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd82;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd82)) begin
            $error("Failed on action=12452 checking port data_out_data. Expected %x, got %x" , 16'd82, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12453 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12454 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12459 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd83;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12464 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12465 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12470 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd84;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd84)) begin
            $error("Failed on action=12475 checking port data_out_data. Expected %x, got %x" , 16'd84, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12476 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12477 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12482 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd85;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12487 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12488 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12493 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd86;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd86)) begin
            $error("Failed on action=12498 checking port data_out_data. Expected %x, got %x" , 16'd86, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12499 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12500 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12505 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd87;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12510 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12511 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd88;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd88)) begin
            $error("Failed on action=12521 checking port data_out_data. Expected %x, got %x" , 16'd88, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12522 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12523 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12528 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd89;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12534 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd90;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd90)) begin
            $error("Failed on action=12544 checking port data_out_data. Expected %x, got %x" , 16'd90, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12545 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12546 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12551 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd91;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12556 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12557 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12562 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd92;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd92)) begin
            $error("Failed on action=12567 checking port data_out_data. Expected %x, got %x" , 16'd92, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12568 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12569 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12574 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd93;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12579 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12580 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12585 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd94;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd94)) begin
            $error("Failed on action=12590 checking port data_out_data. Expected %x, got %x" , 16'd94, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12591 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12592 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12597 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd95;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12602 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12603 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12608 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd96;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12614 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12619 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd97;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12624 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12625 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12630 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd98;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12635 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12636 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12641 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd99;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12646 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12647 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12652 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd100;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12657 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12658 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12663 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd101;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12668 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12669 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12674 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd102;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12679 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12680 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12685 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd103;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12690 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12691 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12696 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd104;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12701 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12702 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12707 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd105;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12712 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12713 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12718 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd106;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12723 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12724 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12729 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd107;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12734 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12735 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12740 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd108;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12745 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12746 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12751 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd109;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12756 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12757 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12762 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd110;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12767 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12768 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12773 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd111;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12779 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12784 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd112;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12789 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12790 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12795 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd113;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12800 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12801 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12806 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd114;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12811 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12812 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12817 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd115;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12822 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12823 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12828 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd116;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12833 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12834 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12839 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd117;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12844 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12845 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12850 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd118;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12855 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12856 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12861 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd119;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12866 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12867 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12872 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd120;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12877 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12878 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12883 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd121;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12888 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12889 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12894 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd122;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12899 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12900 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12905 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd123;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12910 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12911 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd124;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12921 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12922 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12927 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd125;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12932 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12933 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12938 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd126;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12943 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12944 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12949 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd127;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12954 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12955 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12960 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd128;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd128)) begin
            $error("Failed on action=12965 checking port data_out_data. Expected %x, got %x" , 16'd128, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12966 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12967 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12972 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd129;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12977 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12978 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12983 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd130;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd130)) begin
            $error("Failed on action=12988 checking port data_out_data. Expected %x, got %x" , 16'd130, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=12989 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=12990 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=12995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd131;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13000 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13001 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13006 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd132;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd132)) begin
            $error("Failed on action=13011 checking port data_out_data. Expected %x, got %x" , 16'd132, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13012 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13013 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd133;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13023 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13024 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13029 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd134;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd134)) begin
            $error("Failed on action=13034 checking port data_out_data. Expected %x, got %x" , 16'd134, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13035 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13036 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13041 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd135;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13046 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13047 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13052 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd136;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd136)) begin
            $error("Failed on action=13057 checking port data_out_data. Expected %x, got %x" , 16'd136, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13058 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13059 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13064 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd137;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13069 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13070 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13075 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd138;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd138)) begin
            $error("Failed on action=13080 checking port data_out_data. Expected %x, got %x" , 16'd138, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13081 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13082 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13087 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd139;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13092 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13093 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13098 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd140;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd140)) begin
            $error("Failed on action=13103 checking port data_out_data. Expected %x, got %x" , 16'd140, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13104 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13105 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd141;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13116 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd142;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd142)) begin
            $error("Failed on action=13126 checking port data_out_data. Expected %x, got %x" , 16'd142, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13127 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13128 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd143;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13139 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13144 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd144;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd144)) begin
            $error("Failed on action=13149 checking port data_out_data. Expected %x, got %x" , 16'd144, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13150 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13151 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13156 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd145;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13161 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13162 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13167 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd146;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd146)) begin
            $error("Failed on action=13172 checking port data_out_data. Expected %x, got %x" , 16'd146, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13173 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13174 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13179 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd147;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13184 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13185 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13190 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd148;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd148)) begin
            $error("Failed on action=13195 checking port data_out_data. Expected %x, got %x" , 16'd148, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13196 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13197 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13202 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd149;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13207 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13208 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13213 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd150;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd150)) begin
            $error("Failed on action=13218 checking port data_out_data. Expected %x, got %x" , 16'd150, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13219 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13220 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13225 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd151;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13230 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13231 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13236 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd152;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd152)) begin
            $error("Failed on action=13241 checking port data_out_data. Expected %x, got %x" , 16'd152, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13242 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13243 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13248 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd153;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13254 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd154;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd154)) begin
            $error("Failed on action=13264 checking port data_out_data. Expected %x, got %x" , 16'd154, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13265 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13266 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13271 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd155;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13277 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13282 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd156;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd156)) begin
            $error("Failed on action=13287 checking port data_out_data. Expected %x, got %x" , 16'd156, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13288 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13289 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13294 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd157;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13299 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13300 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13305 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd158;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd158)) begin
            $error("Failed on action=13310 checking port data_out_data. Expected %x, got %x" , 16'd158, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13311 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13312 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13317 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd159;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13322 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13323 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13328 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd160;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13333 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13334 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13339 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd161;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13344 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13345 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13350 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd162;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13355 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13356 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13361 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd163;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13366 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13367 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13372 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd164;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13377 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13378 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13383 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd165;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13388 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13389 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13394 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd166;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13399 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13400 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13405 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd167;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13410 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13411 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13416 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd168;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13421 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13422 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13427 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd169;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13432 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13433 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13438 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd170;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13443 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13444 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13449 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd171;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13454 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13455 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13460 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd172;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13465 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13466 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13471 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd173;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13476 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13477 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13482 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd174;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13487 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13488 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13493 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd175;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13499 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13504 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd176;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13509 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13510 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13515 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd177;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13520 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13521 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13526 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd178;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13531 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13532 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13537 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd179;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13542 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13543 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13548 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd180;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13553 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13554 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13559 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd181;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13564 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13565 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13570 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd182;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13575 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13576 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13581 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd183;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13586 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13587 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13592 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd184;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13597 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13598 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13603 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd185;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13608 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13609 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13614 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd186;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13619 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13620 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13625 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd187;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13630 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13631 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd188;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13641 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13642 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13647 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd189;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13652 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13653 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13658 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd190;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13663 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13664 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13669 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd191;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13674 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13675 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13680 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd192;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd192)) begin
            $error("Failed on action=13685 checking port data_out_data. Expected %x, got %x" , 16'd192, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13686 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13687 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd193;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13697 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13698 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13703 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd194;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd194)) begin
            $error("Failed on action=13708 checking port data_out_data. Expected %x, got %x" , 16'd194, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13709 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13710 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd195;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13720 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13721 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13726 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd196;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd196)) begin
            $error("Failed on action=13731 checking port data_out_data. Expected %x, got %x" , 16'd196, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13732 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13733 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13738 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd197;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13743 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13744 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13749 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd198;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd198)) begin
            $error("Failed on action=13754 checking port data_out_data. Expected %x, got %x" , 16'd198, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13755 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13756 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13761 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd199;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13766 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13767 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13772 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd200;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd200)) begin
            $error("Failed on action=13777 checking port data_out_data. Expected %x, got %x" , 16'd200, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13778 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13779 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13784 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd201;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13789 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13790 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13795 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd202;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd202)) begin
            $error("Failed on action=13800 checking port data_out_data. Expected %x, got %x" , 16'd202, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13801 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13802 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13807 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd203;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13812 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13813 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13818 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd204;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd204)) begin
            $error("Failed on action=13823 checking port data_out_data. Expected %x, got %x" , 16'd204, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13824 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13825 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd205;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13836 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd206;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd206)) begin
            $error("Failed on action=13846 checking port data_out_data. Expected %x, got %x" , 16'd206, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13847 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13848 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd207;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13859 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13864 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd208;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd208)) begin
            $error("Failed on action=13869 checking port data_out_data. Expected %x, got %x" , 16'd208, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13870 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13871 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13876 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd209;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13881 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13882 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13887 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd210;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd210)) begin
            $error("Failed on action=13892 checking port data_out_data. Expected %x, got %x" , 16'd210, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13893 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13894 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13899 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd211;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13904 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13905 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13910 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd212;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd212)) begin
            $error("Failed on action=13915 checking port data_out_data. Expected %x, got %x" , 16'd212, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13916 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13917 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13922 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd213;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13927 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13928 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13933 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd214;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd214)) begin
            $error("Failed on action=13938 checking port data_out_data. Expected %x, got %x" , 16'd214, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13939 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13940 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13945 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd215;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13950 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13951 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13956 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd216;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd216)) begin
            $error("Failed on action=13961 checking port data_out_data. Expected %x, got %x" , 16'd216, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13962 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13963 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13968 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd217;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13974 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd218;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd218)) begin
            $error("Failed on action=13984 checking port data_out_data. Expected %x, got %x" , 16'd218, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=13985 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13986 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13991 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd219;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=13996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=13997 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14002 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd220;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd220)) begin
            $error("Failed on action=14007 checking port data_out_data. Expected %x, got %x" , 16'd220, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14008 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14009 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14014 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd221;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14019 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14020 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14025 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd222;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd222)) begin
            $error("Failed on action=14030 checking port data_out_data. Expected %x, got %x" , 16'd222, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14031 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14032 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14037 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd223;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14042 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14043 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14048 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd224;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14053 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14054 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14059 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd225;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14064 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14065 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14070 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd226;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14075 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14076 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14081 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd227;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14086 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14087 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14092 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd228;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14097 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14098 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14103 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd229;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14108 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14109 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14114 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd230;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14119 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14120 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14125 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd231;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14130 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14131 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14136 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd232;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14141 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14142 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14147 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd233;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14152 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14153 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14158 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd234;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14163 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14164 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14169 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd235;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14174 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14175 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14180 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd236;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14185 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14186 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14191 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd237;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14197 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14202 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd238;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14207 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14208 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14213 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd239;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14218 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14219 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14224 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd240;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14229 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14230 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14235 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd241;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14240 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14241 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14246 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd242;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14251 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14252 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14257 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd243;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14262 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14263 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14268 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd244;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14273 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14274 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14279 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd245;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14284 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14285 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14290 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd246;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14295 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14296 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14301 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd247;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14306 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14307 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14312 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd248;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14317 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14318 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14323 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd249;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14328 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14329 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14334 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd250;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14339 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14340 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14345 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd251;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14350 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14351 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14356 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd252;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14361 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14362 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14367 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd253;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14372 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14373 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14378 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd254;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14383 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14384 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14389 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd255;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14394 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14395 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14400 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd256;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd256)) begin
            $error("Failed on action=14405 checking port data_out_data. Expected %x, got %x" , 16'd256, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14406 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14407 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd257;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14417 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14418 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14423 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd258;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd258)) begin
            $error("Failed on action=14428 checking port data_out_data. Expected %x, got %x" , 16'd258, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14429 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14430 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd259;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14440 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14441 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14446 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd260;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd260)) begin
            $error("Failed on action=14451 checking port data_out_data. Expected %x, got %x" , 16'd260, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14452 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14453 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14458 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd261;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14463 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14464 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14469 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd262;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd262)) begin
            $error("Failed on action=14474 checking port data_out_data. Expected %x, got %x" , 16'd262, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14475 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14476 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14481 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd263;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14486 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14487 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14492 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd264;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd264)) begin
            $error("Failed on action=14497 checking port data_out_data. Expected %x, got %x" , 16'd264, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14498 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14499 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14504 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd265;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14509 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14510 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14515 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd266;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd266)) begin
            $error("Failed on action=14520 checking port data_out_data. Expected %x, got %x" , 16'd266, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14521 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14522 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd267;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14532 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14533 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14538 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd268;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd268)) begin
            $error("Failed on action=14543 checking port data_out_data. Expected %x, got %x" , 16'd268, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14544 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14545 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd269;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14556 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd270;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd270)) begin
            $error("Failed on action=14566 checking port data_out_data. Expected %x, got %x" , 16'd270, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14567 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14568 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14573 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd271;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14579 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14584 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd272;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd272)) begin
            $error("Failed on action=14589 checking port data_out_data. Expected %x, got %x" , 16'd272, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14590 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14591 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14596 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd273;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14601 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14602 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14607 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd274;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd274)) begin
            $error("Failed on action=14612 checking port data_out_data. Expected %x, got %x" , 16'd274, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14613 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14614 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14619 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd275;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14624 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14625 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14630 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd276;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd276)) begin
            $error("Failed on action=14635 checking port data_out_data. Expected %x, got %x" , 16'd276, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14636 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14637 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14642 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd277;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14647 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14648 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14653 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd278;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd278)) begin
            $error("Failed on action=14658 checking port data_out_data. Expected %x, got %x" , 16'd278, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14659 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14660 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd279;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14671 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd280;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd280)) begin
            $error("Failed on action=14681 checking port data_out_data. Expected %x, got %x" , 16'd280, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14682 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14683 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14688 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd281;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14694 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14699 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd282;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd282)) begin
            $error("Failed on action=14704 checking port data_out_data. Expected %x, got %x" , 16'd282, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14705 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14706 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14711 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd283;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14716 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14717 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14722 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd284;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd284)) begin
            $error("Failed on action=14727 checking port data_out_data. Expected %x, got %x" , 16'd284, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14728 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14729 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14734 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd285;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14739 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14740 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14745 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd286;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd286)) begin
            $error("Failed on action=14750 checking port data_out_data. Expected %x, got %x" , 16'd286, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=14751 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14752 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14757 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd287;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14762 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14763 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14768 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd288;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14773 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14774 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14779 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd289;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14784 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14785 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14790 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd290;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14795 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14796 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd291;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14806 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14807 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14812 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd292;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14817 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14818 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14823 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd293;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14828 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14829 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14834 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd294;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14839 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14840 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14845 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd295;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14850 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14851 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14856 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd296;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14861 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14862 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14867 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd297;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14872 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14873 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14878 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd298;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14883 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14884 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14889 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd299;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14894 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14895 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14900 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd300;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14905 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14906 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14911 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd301;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14917 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14922 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd302;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14927 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14928 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14933 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd303;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14938 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14939 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14944 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd304;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14949 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14950 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14955 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd305;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14960 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14961 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14966 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd306;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14971 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14972 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14977 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd307;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14982 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14983 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14988 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd308;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14993 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=14994 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=14999 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd309;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15004 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15005 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15010 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd310;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15015 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15016 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15021 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd311;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15026 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15027 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15032 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd312;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15037 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15038 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15043 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd313;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15048 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15049 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15054 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd314;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15059 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15060 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15065 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd315;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15070 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15071 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15076 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd316;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15081 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15082 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15087 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd317;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15092 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15093 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15098 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd318;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15103 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15104 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15109 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd319;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15114 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15115 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15120 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd320;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd320)) begin
            $error("Failed on action=15125 checking port data_out_data. Expected %x, got %x" , 16'd320, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15126 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15127 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd321;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15137 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15138 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15143 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd322;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd322)) begin
            $error("Failed on action=15148 checking port data_out_data. Expected %x, got %x" , 16'd322, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15149 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15150 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd323;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15160 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15161 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15166 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd324;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd324)) begin
            $error("Failed on action=15171 checking port data_out_data. Expected %x, got %x" , 16'd324, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15172 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15173 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15178 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd325;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15183 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15184 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15189 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd326;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd326)) begin
            $error("Failed on action=15194 checking port data_out_data. Expected %x, got %x" , 16'd326, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15195 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15196 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15201 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd327;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15206 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15207 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15212 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd328;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd328)) begin
            $error("Failed on action=15217 checking port data_out_data. Expected %x, got %x" , 16'd328, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15218 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15219 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15224 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd329;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15229 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15230 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15235 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd330;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd330)) begin
            $error("Failed on action=15240 checking port data_out_data. Expected %x, got %x" , 16'd330, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15241 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15242 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd331;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15252 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15253 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15258 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd332;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd332)) begin
            $error("Failed on action=15263 checking port data_out_data. Expected %x, got %x" , 16'd332, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15264 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15265 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd333;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15276 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd334;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd334)) begin
            $error("Failed on action=15286 checking port data_out_data. Expected %x, got %x" , 16'd334, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15287 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15288 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15293 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd335;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15299 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15304 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd336;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd336)) begin
            $error("Failed on action=15309 checking port data_out_data. Expected %x, got %x" , 16'd336, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15310 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15311 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15316 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd337;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15321 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15322 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15327 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd338;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd338)) begin
            $error("Failed on action=15332 checking port data_out_data. Expected %x, got %x" , 16'd338, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15333 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15334 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15339 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd339;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15344 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15345 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15350 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd340;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd340)) begin
            $error("Failed on action=15355 checking port data_out_data. Expected %x, got %x" , 16'd340, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15356 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15357 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15362 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd341;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15367 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15368 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15373 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd342;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd342)) begin
            $error("Failed on action=15378 checking port data_out_data. Expected %x, got %x" , 16'd342, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15379 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15380 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15385 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd343;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15391 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd344;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd344)) begin
            $error("Failed on action=15401 checking port data_out_data. Expected %x, got %x" , 16'd344, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15402 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15403 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15408 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd345;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15414 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15419 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd346;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd346)) begin
            $error("Failed on action=15424 checking port data_out_data. Expected %x, got %x" , 16'd346, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15425 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15426 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15431 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd347;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15436 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15437 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15442 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd348;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd348)) begin
            $error("Failed on action=15447 checking port data_out_data. Expected %x, got %x" , 16'd348, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15448 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15449 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15454 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd349;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15459 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15460 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15465 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd350;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd350)) begin
            $error("Failed on action=15470 checking port data_out_data. Expected %x, got %x" , 16'd350, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15471 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15472 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15477 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd351;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15482 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15483 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15488 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd352;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15493 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15494 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15499 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd353;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15504 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15505 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15510 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd354;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15515 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15516 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd355;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15526 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15527 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15532 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd356;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15537 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15538 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15543 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd357;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15548 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15549 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15554 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd358;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15559 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15560 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15565 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd359;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15570 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15571 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15576 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd360;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15581 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15582 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15587 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd361;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15592 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15593 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15598 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd362;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15603 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15604 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15609 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd363;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15614 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15615 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15620 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd364;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15625 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15626 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15631 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd365;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15637 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15642 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd366;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15647 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15648 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15653 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd367;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15658 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15659 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15664 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd368;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15669 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15670 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15675 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd369;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15680 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15681 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15686 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd370;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15691 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15692 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15697 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd371;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15702 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15703 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15708 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd372;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15713 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15714 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15719 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd373;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15724 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15725 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15730 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd374;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15735 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15736 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15741 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd375;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15746 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15747 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15752 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd376;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15757 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15758 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15763 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd377;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15768 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15769 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15774 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd378;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15779 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15780 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15785 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd379;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15790 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15791 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15796 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd380;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15802 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15807 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd381;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15812 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15813 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15818 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd382;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15823 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15824 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15829 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd383;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15834 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15835 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15840 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd384;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd384)) begin
            $error("Failed on action=15845 checking port data_out_data. Expected %x, got %x" , 16'd384, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15846 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15847 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd385;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15857 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15858 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15863 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd386;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd386)) begin
            $error("Failed on action=15868 checking port data_out_data. Expected %x, got %x" , 16'd386, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15869 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15870 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd387;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15880 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15881 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15886 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd388;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd388)) begin
            $error("Failed on action=15891 checking port data_out_data. Expected %x, got %x" , 16'd388, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15892 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15893 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15898 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd389;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15903 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15904 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15909 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd390;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd390)) begin
            $error("Failed on action=15914 checking port data_out_data. Expected %x, got %x" , 16'd390, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15915 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15916 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15921 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd391;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15926 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15927 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15932 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd392;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd392)) begin
            $error("Failed on action=15937 checking port data_out_data. Expected %x, got %x" , 16'd392, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15938 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15939 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15944 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd393;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15949 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15950 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15955 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd394;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd394)) begin
            $error("Failed on action=15960 checking port data_out_data. Expected %x, got %x" , 16'd394, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15961 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15962 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd395;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15972 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15973 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15978 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd396;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd396)) begin
            $error("Failed on action=15983 checking port data_out_data. Expected %x, got %x" , 16'd396, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=15984 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15985 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd397;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=15995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=15996 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd398;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd398)) begin
            $error("Failed on action=16006 checking port data_out_data. Expected %x, got %x" , 16'd398, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16007 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16008 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16013 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd399;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16019 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16024 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd400;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd400)) begin
            $error("Failed on action=16029 checking port data_out_data. Expected %x, got %x" , 16'd400, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16030 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16031 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16036 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd401;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16041 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16042 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16047 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd402;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd402)) begin
            $error("Failed on action=16052 checking port data_out_data. Expected %x, got %x" , 16'd402, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16053 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16054 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16059 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd403;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16064 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16065 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16070 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd404;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd404)) begin
            $error("Failed on action=16075 checking port data_out_data. Expected %x, got %x" , 16'd404, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16076 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16077 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16082 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd405;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16087 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16088 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16093 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd406;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd406)) begin
            $error("Failed on action=16098 checking port data_out_data. Expected %x, got %x" , 16'd406, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16099 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16100 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16105 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd407;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16111 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd408;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd408)) begin
            $error("Failed on action=16121 checking port data_out_data. Expected %x, got %x" , 16'd408, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16122 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16123 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16128 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd409;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16134 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16139 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd410;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd410)) begin
            $error("Failed on action=16144 checking port data_out_data. Expected %x, got %x" , 16'd410, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16145 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16146 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16151 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd411;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16156 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16157 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16162 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd412;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd412)) begin
            $error("Failed on action=16167 checking port data_out_data. Expected %x, got %x" , 16'd412, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16168 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16169 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16174 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd413;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16179 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16180 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16185 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd414;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd414)) begin
            $error("Failed on action=16190 checking port data_out_data. Expected %x, got %x" , 16'd414, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16191 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16192 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16197 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd415;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16202 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16203 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16208 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd416;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16213 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16214 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd417;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16224 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16225 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16230 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd418;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16235 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16236 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16241 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd419;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16246 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16247 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16252 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd420;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16257 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16258 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16263 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd421;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16268 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16269 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16274 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd422;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16279 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16280 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16285 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd423;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16290 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16291 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16296 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd424;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16301 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16302 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16307 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd425;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16312 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16313 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16318 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd426;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16323 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16324 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16329 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd427;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16334 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16335 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16340 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd428;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16345 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16346 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16351 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd429;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16356 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16357 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16362 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd430;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16367 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16368 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16373 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd431;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16378 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16379 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd432;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16389 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16390 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16395 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd433;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16400 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16401 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16406 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd434;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16411 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16412 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16417 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd435;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16422 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16423 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16428 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd436;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16433 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16434 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16439 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd437;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16444 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16445 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16450 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd438;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16455 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16456 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16461 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd439;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16466 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16467 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16472 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd440;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16477 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16478 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16483 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd441;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16488 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16489 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16494 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd442;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16499 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16500 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16505 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd443;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16510 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16511 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd444;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16522 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd445;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16532 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16533 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16538 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd446;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16543 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16544 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16549 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd447;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16554 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16555 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16560 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd448;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd448)) begin
            $error("Failed on action=16565 checking port data_out_data. Expected %x, got %x" , 16'd448, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16566 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16567 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd449;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16577 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16578 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16583 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd450;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd450)) begin
            $error("Failed on action=16588 checking port data_out_data. Expected %x, got %x" , 16'd450, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16589 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16590 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16595 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd451;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16600 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16601 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16606 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd452;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd452)) begin
            $error("Failed on action=16611 checking port data_out_data. Expected %x, got %x" , 16'd452, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16612 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16613 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16618 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd453;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16623 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16624 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16629 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd454;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd454)) begin
            $error("Failed on action=16634 checking port data_out_data. Expected %x, got %x" , 16'd454, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16635 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16636 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16641 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd455;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16646 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16647 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16652 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd456;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd456)) begin
            $error("Failed on action=16657 checking port data_out_data. Expected %x, got %x" , 16'd456, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16658 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16659 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16664 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd457;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16669 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16670 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16675 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd458;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd458)) begin
            $error("Failed on action=16680 checking port data_out_data. Expected %x, got %x" , 16'd458, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16681 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16682 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd459;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16693 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd460;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd460)) begin
            $error("Failed on action=16703 checking port data_out_data. Expected %x, got %x" , 16'd460, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16704 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16705 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd461;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16716 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16721 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd462;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd462)) begin
            $error("Failed on action=16726 checking port data_out_data. Expected %x, got %x" , 16'd462, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16727 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16728 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16733 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd463;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16738 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16739 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16744 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd464;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd464)) begin
            $error("Failed on action=16749 checking port data_out_data. Expected %x, got %x" , 16'd464, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16750 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16751 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16756 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd465;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16761 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16762 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16767 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd466;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd466)) begin
            $error("Failed on action=16772 checking port data_out_data. Expected %x, got %x" , 16'd466, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16773 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16774 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16779 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd467;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16784 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16785 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16790 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd468;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd468)) begin
            $error("Failed on action=16795 checking port data_out_data. Expected %x, got %x" , 16'd468, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16796 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16797 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16802 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd469;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16807 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16808 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16813 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd470;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd470)) begin
            $error("Failed on action=16818 checking port data_out_data. Expected %x, got %x" , 16'd470, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16819 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16820 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16825 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd471;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16831 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd472;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd472)) begin
            $error("Failed on action=16841 checking port data_out_data. Expected %x, got %x" , 16'd472, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16842 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16843 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16848 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd473;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16854 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16859 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd474;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd474)) begin
            $error("Failed on action=16864 checking port data_out_data. Expected %x, got %x" , 16'd474, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16865 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16866 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16871 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd475;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16876 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16877 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16882 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd476;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd476)) begin
            $error("Failed on action=16887 checking port data_out_data. Expected %x, got %x" , 16'd476, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16888 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16889 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16894 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd477;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16899 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16900 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16905 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd478;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd478)) begin
            $error("Failed on action=16910 checking port data_out_data. Expected %x, got %x" , 16'd478, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=16911 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16912 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16917 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd479;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16922 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16923 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16928 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd480;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16933 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16934 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd481;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16944 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16945 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16950 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd482;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16955 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16956 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16961 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd483;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16966 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16967 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16972 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd484;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16977 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16978 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16983 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd485;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16988 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=16989 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16994 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd486;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=16999 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17000 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17005 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd487;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17010 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17011 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17016 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd488;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17021 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17022 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17027 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd489;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17032 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17033 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17038 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd490;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17043 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17044 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17049 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd491;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17054 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17055 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17060 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd492;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17065 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17066 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17071 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd493;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17076 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17077 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17082 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd494;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17087 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17088 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17093 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd495;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17098 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17099 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd496;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17109 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17110 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd497;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17120 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17121 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17126 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd498;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17131 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17132 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17137 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd499;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17142 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17143 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17148 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd500;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17153 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17154 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17159 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd501;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17164 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17165 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17170 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd502;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17175 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17176 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17181 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd503;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17186 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17187 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17192 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd504;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17197 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17198 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17203 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd505;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17208 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17209 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17214 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd506;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17220 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17225 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd507;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17230 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17231 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17236 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd508;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17241 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17242 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd509;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17252 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17253 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17258 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd510;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17263 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17264 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17269 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd511;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17274 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17275 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17280 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd512;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd512)) begin
            $error("Failed on action=17285 checking port data_out_data. Expected %x, got %x" , 16'd512, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17286 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17287 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd513;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17297 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17298 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17303 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd514;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd514)) begin
            $error("Failed on action=17308 checking port data_out_data. Expected %x, got %x" , 16'd514, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17309 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17310 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17315 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd515;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17320 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17321 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17326 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd516;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd516)) begin
            $error("Failed on action=17331 checking port data_out_data. Expected %x, got %x" , 16'd516, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17332 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17333 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17338 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd517;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17343 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17344 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17349 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd518;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd518)) begin
            $error("Failed on action=17354 checking port data_out_data. Expected %x, got %x" , 16'd518, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17355 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17356 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17361 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd519;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17366 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17367 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17372 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd520;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd520)) begin
            $error("Failed on action=17377 checking port data_out_data. Expected %x, got %x" , 16'd520, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17378 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17379 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd521;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17389 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17390 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17395 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd522;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd522)) begin
            $error("Failed on action=17400 checking port data_out_data. Expected %x, got %x" , 16'd522, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17401 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17402 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd523;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17413 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd524;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd524)) begin
            $error("Failed on action=17423 checking port data_out_data. Expected %x, got %x" , 16'd524, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17424 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17425 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17430 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd525;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17436 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17441 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd526;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd526)) begin
            $error("Failed on action=17446 checking port data_out_data. Expected %x, got %x" , 16'd526, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17447 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17448 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17453 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd527;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17458 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17459 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17464 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd528;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd528)) begin
            $error("Failed on action=17469 checking port data_out_data. Expected %x, got %x" , 16'd528, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17470 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17471 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17476 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd529;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17481 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17482 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17487 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd530;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd530)) begin
            $error("Failed on action=17492 checking port data_out_data. Expected %x, got %x" , 16'd530, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17493 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17494 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17499 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd531;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17504 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17505 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17510 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd532;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd532)) begin
            $error("Failed on action=17515 checking port data_out_data. Expected %x, got %x" , 16'd532, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17516 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17517 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17522 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd533;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17528 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd534;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd534)) begin
            $error("Failed on action=17538 checking port data_out_data. Expected %x, got %x" , 16'd534, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17539 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17540 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17545 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd535;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17551 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17556 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd536;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd536)) begin
            $error("Failed on action=17561 checking port data_out_data. Expected %x, got %x" , 16'd536, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17562 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17563 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17568 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd537;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17573 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17574 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17579 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd538;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd538)) begin
            $error("Failed on action=17584 checking port data_out_data. Expected %x, got %x" , 16'd538, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17585 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17586 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17591 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd539;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17596 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17597 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17602 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd540;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd540)) begin
            $error("Failed on action=17607 checking port data_out_data. Expected %x, got %x" , 16'd540, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17608 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17609 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17614 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd541;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17619 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17620 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17625 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd542;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd542)) begin
            $error("Failed on action=17630 checking port data_out_data. Expected %x, got %x" , 16'd542, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=17631 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17632 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17637 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd543;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17642 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17643 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17648 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd544;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17653 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17654 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd545;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17664 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17665 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd546;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17675 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17676 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd547;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17686 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17687 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd548;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17697 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17698 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17703 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd549;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17708 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17709 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17714 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd550;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17719 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17720 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17725 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd551;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17730 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17731 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17736 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd552;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17741 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17742 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17747 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd553;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17752 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17753 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17758 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd554;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17763 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17764 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17769 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd555;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17774 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17775 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17780 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd556;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17785 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17786 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17791 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd557;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17796 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17797 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17802 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd558;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17807 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17808 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17813 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd559;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17818 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17819 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd560;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17829 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17830 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd561;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17840 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17841 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17846 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd562;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17851 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17852 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17857 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd563;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17862 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17863 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17868 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd564;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17873 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17874 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17879 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd565;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17884 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17885 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17890 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd566;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17895 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17896 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17901 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd567;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17906 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17907 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17912 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd568;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17917 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17918 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17923 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd569;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17928 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17929 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17934 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd570;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17940 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17945 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd571;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17950 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17951 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17956 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd572;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17961 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17962 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd573;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17972 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17973 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17978 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd574;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17983 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17984 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17989 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd575;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=17994 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=17995 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18000 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd576;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd576)) begin
            $error("Failed on action=18005 checking port data_out_data. Expected %x, got %x" , 16'd576, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18006 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18007 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd577;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18017 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18018 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18023 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd578;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd578)) begin
            $error("Failed on action=18028 checking port data_out_data. Expected %x, got %x" , 16'd578, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18029 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18030 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18035 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd579;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18040 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18041 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18046 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd580;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd580)) begin
            $error("Failed on action=18051 checking port data_out_data. Expected %x, got %x" , 16'd580, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18052 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18053 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18058 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd581;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18063 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18064 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18069 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd582;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd582)) begin
            $error("Failed on action=18074 checking port data_out_data. Expected %x, got %x" , 16'd582, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18075 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18076 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18081 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd583;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18086 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18087 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18092 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd584;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd584)) begin
            $error("Failed on action=18097 checking port data_out_data. Expected %x, got %x" , 16'd584, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18098 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18099 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd585;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18109 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18110 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd586;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd586)) begin
            $error("Failed on action=18120 checking port data_out_data. Expected %x, got %x" , 16'd586, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18121 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18122 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd587;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18133 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd588;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd588)) begin
            $error("Failed on action=18143 checking port data_out_data. Expected %x, got %x" , 16'd588, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18144 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18145 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd589;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18156 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18161 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd590;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd590)) begin
            $error("Failed on action=18166 checking port data_out_data. Expected %x, got %x" , 16'd590, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18167 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18168 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd591;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18178 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18179 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18184 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd592;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd592)) begin
            $error("Failed on action=18189 checking port data_out_data. Expected %x, got %x" , 16'd592, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18190 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18191 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd593;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18201 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18202 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18207 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd594;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd594)) begin
            $error("Failed on action=18212 checking port data_out_data. Expected %x, got %x" , 16'd594, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18213 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18214 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd595;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18224 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18225 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18230 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd596;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd596)) begin
            $error("Failed on action=18235 checking port data_out_data. Expected %x, got %x" , 16'd596, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18236 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18237 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd597;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18248 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd598;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd598)) begin
            $error("Failed on action=18258 checking port data_out_data. Expected %x, got %x" , 16'd598, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18259 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18260 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18265 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd599;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18271 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd600;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd600)) begin
            $error("Failed on action=18281 checking port data_out_data. Expected %x, got %x" , 16'd600, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18282 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18283 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18288 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd601;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18293 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18294 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18299 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd602;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd602)) begin
            $error("Failed on action=18304 checking port data_out_data. Expected %x, got %x" , 16'd602, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18305 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18306 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18311 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd603;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18316 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18317 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18322 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd604;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd604)) begin
            $error("Failed on action=18327 checking port data_out_data. Expected %x, got %x" , 16'd604, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18328 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18329 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18334 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd605;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18339 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18340 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18345 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd606;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd606)) begin
            $error("Failed on action=18350 checking port data_out_data. Expected %x, got %x" , 16'd606, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18351 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18352 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18357 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd607;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18362 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18363 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18368 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd608;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18373 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18374 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd609;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18385 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd610;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18395 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18396 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd611;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18406 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18407 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd612;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18417 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18418 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18423 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd613;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18428 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18429 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18434 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd614;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18439 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18440 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18445 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd615;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18450 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18451 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18456 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd616;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18461 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18462 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18467 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd617;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18472 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18473 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18478 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd618;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18483 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18484 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18489 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd619;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18494 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18495 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18500 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd620;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18505 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18506 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18511 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd621;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18517 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18522 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd622;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18528 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd623;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18538 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18539 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd624;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18549 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18550 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd625;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18560 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18561 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18566 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd626;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18571 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18572 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18577 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd627;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18582 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18583 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18588 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd628;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18593 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18594 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18599 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd629;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18604 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18605 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18610 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd630;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18615 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18616 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18621 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd631;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18626 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18627 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18632 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd632;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18637 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18638 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18643 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd633;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18648 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18649 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18654 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd634;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18660 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd635;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18671 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd636;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18682 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd637;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18693 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd638;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18703 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18704 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd639;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18714 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18715 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18720 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd640;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd640)) begin
            $error("Failed on action=18725 checking port data_out_data. Expected %x, got %x" , 16'd640, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18726 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18727 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd641;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18737 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18738 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18743 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd642;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd642)) begin
            $error("Failed on action=18748 checking port data_out_data. Expected %x, got %x" , 16'd642, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18749 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18750 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd643;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18760 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18761 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18766 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd644;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd644)) begin
            $error("Failed on action=18771 checking port data_out_data. Expected %x, got %x" , 16'd644, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18772 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18773 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd645;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18783 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18784 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18789 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd646;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd646)) begin
            $error("Failed on action=18794 checking port data_out_data. Expected %x, got %x" , 16'd646, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18795 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18796 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd647;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18806 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18807 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18812 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd648;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd648)) begin
            $error("Failed on action=18817 checking port data_out_data. Expected %x, got %x" , 16'd648, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18818 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18819 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd649;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18829 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18830 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd650;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd650)) begin
            $error("Failed on action=18840 checking port data_out_data. Expected %x, got %x" , 16'd650, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18841 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18842 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd651;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18853 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd652;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd652)) begin
            $error("Failed on action=18863 checking port data_out_data. Expected %x, got %x" , 16'd652, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18864 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18865 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd653;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18876 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18881 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd654;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd654)) begin
            $error("Failed on action=18886 checking port data_out_data. Expected %x, got %x" , 16'd654, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18887 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18888 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd655;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18898 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18899 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18904 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd656;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd656)) begin
            $error("Failed on action=18909 checking port data_out_data. Expected %x, got %x" , 16'd656, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18910 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18911 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd657;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18921 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18922 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18927 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd658;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd658)) begin
            $error("Failed on action=18932 checking port data_out_data. Expected %x, got %x" , 16'd658, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18933 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18934 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd659;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18944 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18945 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18950 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd660;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd660)) begin
            $error("Failed on action=18955 checking port data_out_data. Expected %x, got %x" , 16'd660, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18956 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18957 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd661;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18968 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd662;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd662)) begin
            $error("Failed on action=18978 checking port data_out_data. Expected %x, got %x" , 16'd662, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=18979 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18980 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18985 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd663;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=18991 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=18996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd664;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd664)) begin
            $error("Failed on action=19001 checking port data_out_data. Expected %x, got %x" , 16'd664, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19002 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19003 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19008 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd665;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19013 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19014 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19019 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd666;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd666)) begin
            $error("Failed on action=19024 checking port data_out_data. Expected %x, got %x" , 16'd666, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19025 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19026 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19031 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd667;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19036 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19037 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19042 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd668;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd668)) begin
            $error("Failed on action=19047 checking port data_out_data. Expected %x, got %x" , 16'd668, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19048 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19049 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19054 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd669;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19059 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19060 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19065 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd670;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd670)) begin
            $error("Failed on action=19070 checking port data_out_data. Expected %x, got %x" , 16'd670, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19071 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19072 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19077 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd671;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19082 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19083 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19088 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd672;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19093 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19094 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd673;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19105 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd674;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19115 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19116 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd675;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19126 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19127 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd676;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19137 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19138 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19143 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd677;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19148 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19149 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19154 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd678;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19159 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19160 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19165 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd679;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19170 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19171 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19176 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd680;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19181 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19182 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19187 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd681;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19192 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19193 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19198 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd682;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19203 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19204 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19209 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd683;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19214 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19215 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19220 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd684;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19225 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19226 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19231 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd685;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19236 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19237 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd686;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19247 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19248 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd687;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19258 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19259 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd688;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19269 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19270 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd689;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19280 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19281 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19286 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd690;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19291 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19292 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19297 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd691;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19302 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19303 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19308 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd692;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19313 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19314 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19319 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd693;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19324 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19325 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19330 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd694;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19335 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19336 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19341 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd695;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19346 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19347 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19352 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd696;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19357 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19358 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19363 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd697;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19368 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19369 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19374 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd698;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19380 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19385 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd699;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19391 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd700;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19402 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd701;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19413 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd702;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19423 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19424 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd703;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19434 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19435 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19440 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd704;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd704)) begin
            $error("Failed on action=19445 checking port data_out_data. Expected %x, got %x" , 16'd704, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19446 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19447 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd705;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19457 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19458 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19463 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd706;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd706)) begin
            $error("Failed on action=19468 checking port data_out_data. Expected %x, got %x" , 16'd706, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19469 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19470 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd707;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19480 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19481 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19486 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd708;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd708)) begin
            $error("Failed on action=19491 checking port data_out_data. Expected %x, got %x" , 16'd708, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19492 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19493 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd709;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19503 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19504 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19509 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd710;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd710)) begin
            $error("Failed on action=19514 checking port data_out_data. Expected %x, got %x" , 16'd710, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19515 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19516 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd711;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19526 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19527 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19532 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd712;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd712)) begin
            $error("Failed on action=19537 checking port data_out_data. Expected %x, got %x" , 16'd712, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19538 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19539 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd713;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19549 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19550 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd714;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd714)) begin
            $error("Failed on action=19560 checking port data_out_data. Expected %x, got %x" , 16'd714, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19561 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19562 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd715;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19573 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd716;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd716)) begin
            $error("Failed on action=19583 checking port data_out_data. Expected %x, got %x" , 16'd716, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19584 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19585 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd717;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19595 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19596 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19601 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd718;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd718)) begin
            $error("Failed on action=19606 checking port data_out_data. Expected %x, got %x" , 16'd718, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19607 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19608 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd719;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19618 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19619 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19624 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd720;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd720)) begin
            $error("Failed on action=19629 checking port data_out_data. Expected %x, got %x" , 16'd720, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19630 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19631 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd721;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19641 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19642 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19647 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd722;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd722)) begin
            $error("Failed on action=19652 checking port data_out_data. Expected %x, got %x" , 16'd722, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19653 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19654 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd723;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19664 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19665 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19670 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd724;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd724)) begin
            $error("Failed on action=19675 checking port data_out_data. Expected %x, got %x" , 16'd724, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19676 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19677 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd725;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19688 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd726;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd726)) begin
            $error("Failed on action=19698 checking port data_out_data. Expected %x, got %x" , 16'd726, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19699 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19700 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19705 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd727;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19711 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19716 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd728;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd728)) begin
            $error("Failed on action=19721 checking port data_out_data. Expected %x, got %x" , 16'd728, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19722 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19723 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19728 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd729;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19733 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19734 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19739 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd730;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd730)) begin
            $error("Failed on action=19744 checking port data_out_data. Expected %x, got %x" , 16'd730, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19745 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19746 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19751 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd731;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19756 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19757 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19762 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd732;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd732)) begin
            $error("Failed on action=19767 checking port data_out_data. Expected %x, got %x" , 16'd732, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19768 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19769 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19774 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd733;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19779 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19780 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19785 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd734;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd734)) begin
            $error("Failed on action=19790 checking port data_out_data. Expected %x, got %x" , 16'd734, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=19791 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19792 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19797 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd735;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19802 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19803 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19808 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd736;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19813 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19814 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd737;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19825 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd738;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19835 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19836 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd739;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19846 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19847 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd740;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19857 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19858 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19863 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd741;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19868 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19869 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19874 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd742;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19879 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19880 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19885 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd743;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19890 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19891 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19896 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd744;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19901 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19902 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19907 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd745;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19912 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19913 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19918 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd746;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19923 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19924 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19929 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd747;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19934 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19935 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19940 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd748;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19945 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19946 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19951 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd749;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19956 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19957 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd750;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19967 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19968 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd751;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19978 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19979 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd752;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19989 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=19990 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=19995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd753;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20000 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20001 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20006 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd754;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20011 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20012 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20017 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd755;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20022 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20023 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20028 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd756;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20033 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20034 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20039 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd757;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20044 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20045 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20050 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd758;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20055 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20056 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20061 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd759;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20066 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20067 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20072 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd760;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20077 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20078 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20083 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd761;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20088 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20089 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20094 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd762;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20100 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20105 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd763;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20111 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd764;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20121 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20122 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd765;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20132 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20133 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd766;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20143 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20144 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20149 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd767;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20154 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20155 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20160 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd768;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd768)) begin
            $error("Failed on action=20165 checking port data_out_data. Expected %x, got %x" , 16'd768, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20166 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20167 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20172 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd769;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20177 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20178 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20183 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd770;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd770)) begin
            $error("Failed on action=20188 checking port data_out_data. Expected %x, got %x" , 16'd770, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20189 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20190 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20195 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd771;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20200 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20201 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20206 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd772;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd772)) begin
            $error("Failed on action=20211 checking port data_out_data. Expected %x, got %x" , 16'd772, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20212 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20213 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20218 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd773;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20223 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20224 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20229 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd774;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd774)) begin
            $error("Failed on action=20234 checking port data_out_data. Expected %x, got %x" , 16'd774, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20235 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20236 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20241 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd775;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20246 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20247 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20252 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd776;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd776)) begin
            $error("Failed on action=20257 checking port data_out_data. Expected %x, got %x" , 16'd776, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20258 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20259 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd777;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20269 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20270 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd778;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd778)) begin
            $error("Failed on action=20280 checking port data_out_data. Expected %x, got %x" , 16'd778, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20281 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20282 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd779;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20293 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd780;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd780)) begin
            $error("Failed on action=20303 checking port data_out_data. Expected %x, got %x" , 16'd780, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20304 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20305 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20310 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd781;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20315 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20316 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20321 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd782;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd782)) begin
            $error("Failed on action=20326 checking port data_out_data. Expected %x, got %x" , 16'd782, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20327 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20328 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20333 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd783;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20338 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20339 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20344 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd784;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd784)) begin
            $error("Failed on action=20349 checking port data_out_data. Expected %x, got %x" , 16'd784, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20350 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20351 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20356 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd785;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20361 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20362 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20367 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd786;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd786)) begin
            $error("Failed on action=20372 checking port data_out_data. Expected %x, got %x" , 16'd786, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20373 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20374 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20379 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd787;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20384 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20385 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20390 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd788;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd788)) begin
            $error("Failed on action=20395 checking port data_out_data. Expected %x, got %x" , 16'd788, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20396 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20397 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20402 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd789;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20408 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd790;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd790)) begin
            $error("Failed on action=20418 checking port data_out_data. Expected %x, got %x" , 16'd790, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20419 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20420 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20425 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd791;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20430 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20431 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20436 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd792;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd792)) begin
            $error("Failed on action=20441 checking port data_out_data. Expected %x, got %x" , 16'd792, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20442 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20443 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20448 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd793;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20453 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20454 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20459 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd794;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd794)) begin
            $error("Failed on action=20464 checking port data_out_data. Expected %x, got %x" , 16'd794, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20465 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20466 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20471 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd795;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20476 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20477 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20482 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd796;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd796)) begin
            $error("Failed on action=20487 checking port data_out_data. Expected %x, got %x" , 16'd796, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20488 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20489 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20494 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd797;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20499 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20500 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20505 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd798;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd798)) begin
            $error("Failed on action=20510 checking port data_out_data. Expected %x, got %x" , 16'd798, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20511 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20512 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20517 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd799;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20522 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20523 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20528 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd800;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20533 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20534 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd801;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20545 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd802;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20555 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20556 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd803;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20566 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20567 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd804;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20577 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20578 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20583 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd805;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20588 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20589 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20594 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd806;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20599 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20600 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20605 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd807;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20610 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20611 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20616 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd808;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20621 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20622 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20627 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd809;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20632 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20633 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20638 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd810;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20643 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20644 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20649 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd811;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20654 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20655 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20660 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd812;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20666 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20671 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd813;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20676 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20677 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd814;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20687 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20688 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd815;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20698 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20699 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd816;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20710 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd817;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20720 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20721 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20726 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd818;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20731 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20732 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20737 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd819;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20742 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20743 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20748 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd820;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20753 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20754 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20759 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd821;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20764 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20765 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20770 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd822;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20775 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20776 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20781 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd823;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20786 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20787 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20792 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd824;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20797 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20798 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20803 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd825;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20808 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20809 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20814 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd826;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20820 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20825 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd827;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20831 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd828;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20841 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20842 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd829;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20852 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20853 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd830;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20863 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20864 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20869 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd831;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20874 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20875 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20880 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd832;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd832)) begin
            $error("Failed on action=20885 checking port data_out_data. Expected %x, got %x" , 16'd832, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20886 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20887 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20892 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd833;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20897 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20898 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20903 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd834;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd834)) begin
            $error("Failed on action=20908 checking port data_out_data. Expected %x, got %x" , 16'd834, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20909 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20910 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20915 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd835;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20920 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20921 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20926 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd836;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd836)) begin
            $error("Failed on action=20931 checking port data_out_data. Expected %x, got %x" , 16'd836, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20932 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20933 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20938 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd837;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20943 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20944 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20949 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd838;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd838)) begin
            $error("Failed on action=20954 checking port data_out_data. Expected %x, got %x" , 16'd838, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20955 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20956 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20961 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd839;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20966 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20967 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20972 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd840;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd840)) begin
            $error("Failed on action=20977 checking port data_out_data. Expected %x, got %x" , 16'd840, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=20978 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20979 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd841;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20989 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=20990 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=20995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd842;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd842)) begin
            $error("Failed on action=21000 checking port data_out_data. Expected %x, got %x" , 16'd842, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21001 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21002 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd843;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21013 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd844;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd844)) begin
            $error("Failed on action=21023 checking port data_out_data. Expected %x, got %x" , 16'd844, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21024 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21025 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21030 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd845;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21035 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21036 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21041 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd846;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd846)) begin
            $error("Failed on action=21046 checking port data_out_data. Expected %x, got %x" , 16'd846, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21047 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21048 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21053 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd847;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21058 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21059 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21064 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd848;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd848)) begin
            $error("Failed on action=21069 checking port data_out_data. Expected %x, got %x" , 16'd848, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21070 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21071 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21076 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd849;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21081 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21082 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21087 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd850;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd850)) begin
            $error("Failed on action=21092 checking port data_out_data. Expected %x, got %x" , 16'd850, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21093 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21094 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21099 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd851;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21104 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21105 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21110 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd852;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd852)) begin
            $error("Failed on action=21115 checking port data_out_data. Expected %x, got %x" , 16'd852, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21116 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21117 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21122 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd853;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21128 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd854;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd854)) begin
            $error("Failed on action=21138 checking port data_out_data. Expected %x, got %x" , 16'd854, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21139 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21140 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21145 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd855;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21150 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21151 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21156 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd856;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd856)) begin
            $error("Failed on action=21161 checking port data_out_data. Expected %x, got %x" , 16'd856, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21162 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21163 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21168 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd857;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21173 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21174 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21179 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd858;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd858)) begin
            $error("Failed on action=21184 checking port data_out_data. Expected %x, got %x" , 16'd858, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21185 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21186 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21191 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd859;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21196 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21197 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21202 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd860;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd860)) begin
            $error("Failed on action=21207 checking port data_out_data. Expected %x, got %x" , 16'd860, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21208 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21209 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21214 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd861;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21219 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21220 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21225 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd862;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd862)) begin
            $error("Failed on action=21230 checking port data_out_data. Expected %x, got %x" , 16'd862, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21231 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21232 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21237 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd863;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21242 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21243 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21248 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd864;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21253 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21254 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd865;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21264 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21265 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd866;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21275 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21276 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd867;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21286 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21287 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd868;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21297 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21298 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21303 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd869;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21308 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21309 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21314 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd870;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21319 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21320 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21325 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd871;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21330 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21331 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21336 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd872;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21341 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21342 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21347 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd873;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21352 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21353 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21358 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd874;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21363 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21364 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21369 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd875;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21374 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21375 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21380 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd876;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21385 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21386 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21391 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd877;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21396 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21397 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21402 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd878;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21407 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21408 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21413 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd879;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21418 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21419 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd880;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21430 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd881;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21440 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21441 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21446 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd882;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21451 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21452 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21457 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd883;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21462 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21463 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21468 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd884;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21473 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21474 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21479 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd885;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21484 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21485 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21490 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd886;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21495 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21496 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21501 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd887;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21506 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21507 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21512 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd888;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21517 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21518 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21523 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd889;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21528 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21529 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21534 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd890;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21540 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21545 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd891;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21551 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21556 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd892;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21561 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21562 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd893;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21572 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21573 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21578 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd894;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21583 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21584 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21589 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd895;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21594 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21595 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21600 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd896;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd896)) begin
            $error("Failed on action=21605 checking port data_out_data. Expected %x, got %x" , 16'd896, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21606 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21607 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21612 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd897;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21617 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21618 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21623 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd898;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd898)) begin
            $error("Failed on action=21628 checking port data_out_data. Expected %x, got %x" , 16'd898, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21629 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21630 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21635 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd899;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21640 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21641 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21646 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd900;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd900)) begin
            $error("Failed on action=21651 checking port data_out_data. Expected %x, got %x" , 16'd900, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21652 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21653 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21658 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd901;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21663 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21664 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21669 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd902;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd902)) begin
            $error("Failed on action=21674 checking port data_out_data. Expected %x, got %x" , 16'd902, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21675 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21676 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21681 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd903;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21686 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21687 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21692 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd904;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd904)) begin
            $error("Failed on action=21697 checking port data_out_data. Expected %x, got %x" , 16'd904, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21698 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21699 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd905;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21709 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21710 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd906;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd906)) begin
            $error("Failed on action=21720 checking port data_out_data. Expected %x, got %x" , 16'd906, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21721 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21722 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21727 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd907;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21733 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21738 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd908;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd908)) begin
            $error("Failed on action=21743 checking port data_out_data. Expected %x, got %x" , 16'd908, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21744 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21745 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21750 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd909;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21755 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21756 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21761 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd910;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd910)) begin
            $error("Failed on action=21766 checking port data_out_data. Expected %x, got %x" , 16'd910, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21767 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21768 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21773 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd911;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21778 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21779 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21784 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd912;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd912)) begin
            $error("Failed on action=21789 checking port data_out_data. Expected %x, got %x" , 16'd912, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21790 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21791 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21796 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd913;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21801 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21802 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21807 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd914;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd914)) begin
            $error("Failed on action=21812 checking port data_out_data. Expected %x, got %x" , 16'd914, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21813 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21814 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21819 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd915;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21824 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21825 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21830 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd916;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd916)) begin
            $error("Failed on action=21835 checking port data_out_data. Expected %x, got %x" , 16'd916, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21836 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21837 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21842 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd917;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21848 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd918;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd918)) begin
            $error("Failed on action=21858 checking port data_out_data. Expected %x, got %x" , 16'd918, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21859 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21860 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21865 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd919;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21870 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21871 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21876 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd920;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd920)) begin
            $error("Failed on action=21881 checking port data_out_data. Expected %x, got %x" , 16'd920, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21882 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21883 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21888 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd921;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21893 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21894 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21899 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd922;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd922)) begin
            $error("Failed on action=21904 checking port data_out_data. Expected %x, got %x" , 16'd922, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21905 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21906 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21911 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd923;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21916 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21917 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21922 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd924;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd924)) begin
            $error("Failed on action=21927 checking port data_out_data. Expected %x, got %x" , 16'd924, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21928 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21929 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21934 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd925;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21939 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21940 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21945 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd926;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd926)) begin
            $error("Failed on action=21950 checking port data_out_data. Expected %x, got %x" , 16'd926, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=21951 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21952 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21957 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd927;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21962 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21963 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21968 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd928;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21973 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21974 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd929;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21984 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21985 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd930;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=21995 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=21996 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd931;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22006 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22007 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd932;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22017 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22018 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22023 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd933;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22028 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22029 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22034 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd934;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22039 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22040 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22045 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd935;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22050 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22051 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22056 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd936;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22061 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22062 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22067 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd937;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22072 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22073 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22078 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd938;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22083 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22084 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22089 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd939;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22094 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22095 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22100 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd940;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22105 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22106 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22111 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd941;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22116 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22117 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22122 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd942;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22127 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22128 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22133 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd943;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22138 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22139 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22144 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd944;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22149 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22150 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22155 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd945;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22160 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22161 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22166 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd946;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22171 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22172 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22177 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd947;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22182 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22183 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22188 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd948;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22193 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22194 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22199 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd949;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22204 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22205 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22210 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd950;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22215 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22216 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22221 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd951;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22226 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22227 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22232 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd952;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22237 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22238 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22243 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd953;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22248 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22249 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22254 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd954;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22259 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22260 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22265 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd955;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22270 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22271 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22276 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd956;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22281 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22282 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22287 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd957;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22292 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22293 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22298 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd958;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22303 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22304 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22309 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd959;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22314 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22315 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22320 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd960;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd960)) begin
            $error("Failed on action=22325 checking port data_out_data. Expected %x, got %x" , 16'd960, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22326 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22327 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22332 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd961;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22337 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22338 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22343 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd962;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd962)) begin
            $error("Failed on action=22348 checking port data_out_data. Expected %x, got %x" , 16'd962, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22349 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22350 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22355 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd963;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22360 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22361 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22366 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd964;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd964)) begin
            $error("Failed on action=22371 checking port data_out_data. Expected %x, got %x" , 16'd964, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22372 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22373 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22378 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd965;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22383 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22384 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22389 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd966;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd966)) begin
            $error("Failed on action=22394 checking port data_out_data. Expected %x, got %x" , 16'd966, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22395 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22396 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22401 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd967;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22406 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22407 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22412 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd968;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd968)) begin
            $error("Failed on action=22417 checking port data_out_data. Expected %x, got %x" , 16'd968, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22418 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22419 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22424 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd969;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22429 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22430 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22435 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd970;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd970)) begin
            $error("Failed on action=22440 checking port data_out_data. Expected %x, got %x" , 16'd970, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22441 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22442 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22447 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd971;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22452 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22453 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22458 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd972;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd972)) begin
            $error("Failed on action=22463 checking port data_out_data. Expected %x, got %x" , 16'd972, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22464 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22465 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22470 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd973;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22475 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22476 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22481 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd974;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd974)) begin
            $error("Failed on action=22486 checking port data_out_data. Expected %x, got %x" , 16'd974, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22487 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22488 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22493 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd975;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22498 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22499 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22504 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd976;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd976)) begin
            $error("Failed on action=22509 checking port data_out_data. Expected %x, got %x" , 16'd976, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22510 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22511 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22516 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd977;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22521 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22522 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22527 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd978;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd978)) begin
            $error("Failed on action=22532 checking port data_out_data. Expected %x, got %x" , 16'd978, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22533 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22534 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22539 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd979;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22544 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22545 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22550 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd980;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd980)) begin
            $error("Failed on action=22555 checking port data_out_data. Expected %x, got %x" , 16'd980, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22556 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22557 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22562 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd981;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22567 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22568 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22573 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd982;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd982)) begin
            $error("Failed on action=22578 checking port data_out_data. Expected %x, got %x" , 16'd982, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22579 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22580 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22585 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd983;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22590 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22591 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22596 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd984;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd984)) begin
            $error("Failed on action=22601 checking port data_out_data. Expected %x, got %x" , 16'd984, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22602 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22603 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22608 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd985;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22613 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22614 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22619 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd986;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd986)) begin
            $error("Failed on action=22624 checking port data_out_data. Expected %x, got %x" , 16'd986, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22625 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22626 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22631 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd987;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22636 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22637 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22642 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd988;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd988)) begin
            $error("Failed on action=22647 checking port data_out_data. Expected %x, got %x" , 16'd988, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22648 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22649 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22654 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd989;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22659 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22660 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22665 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd990;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_data == 16'd990)) begin
            $error("Failed on action=22670 checking port data_out_data. Expected %x, got %x" , 16'd990, data_out_data);

        end
        if (!(data_out_valid == 1'd1)) begin
            $error("Failed on action=22671 checking port data_out_valid. Expected %x, got %x" , 1'd1, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22672 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22677 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd991;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22682 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22683 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22688 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd992;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22693 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22694 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22699 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd993;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22704 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22705 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22710 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd994;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22715 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22716 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22721 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd995;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22726 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22727 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22732 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd996;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22737 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22738 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22743 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd997;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22748 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22749 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22754 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd998;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22759 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22760 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22765 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd999;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22770 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22771 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22776 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1000;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22781 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22782 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22787 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1001;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22792 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22793 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22798 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1002;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22803 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22804 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22809 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1003;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22814 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22815 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22820 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1004;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22825 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22826 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22831 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1005;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22836 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22837 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22842 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1006;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22847 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22848 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22853 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1007;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22858 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22859 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22864 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1008;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22869 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22870 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22875 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1009;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22880 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22881 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22886 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1010;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22891 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22892 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22897 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1011;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22902 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22903 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22908 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1012;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22913 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22914 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22919 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1013;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22924 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22925 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22930 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1014;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22935 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22936 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22941 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1015;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22946 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22947 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22952 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1016;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22957 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22958 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22963 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1017;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22968 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22969 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22974 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1018;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22979 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22980 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22985 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1019;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22990 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=22991 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=22996 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1020;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23001 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=23002 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23007 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1021;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23012 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=23013 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23018 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1022;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23023 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=23024 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23029 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        data_in_valid = 1'd1;
        #5;
        data_in_data = 16'd1023;
        #5;
        data_out_ready = 1'd1;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23034 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end
        if (!(data_in_ready == 1'd1)) begin
            $error("Failed on action=23035 checking port data_in_ready. Expected %x, got %x" , 1'd1, data_in_ready);

        end
        #5 CLK ^= 1;
        #5 CLK ^= 1;
        data_in_valid = 1'd0;
        #5;
        data_out_ready = 1'd0;
        #5;
        if (!(data_out_valid == 1'd0)) begin
            $error("Failed on action=23040 checking port data_out_valid. Expected %x, got %x" , 1'd0, data_out_valid);

        end

        #20 $finish;
    end

endmodule
